// Contributed by Jessica Hausman <Jessica.K.Hausman AT jpl DOT nasa DOT gov>

netcdf cyg.ddmi.s20140920-120002-e20140920-134000.l2.v01.v01 {
dimensions:
	sample = 17839 ;
	num_time_avg_ddms = 5 ;
variables:
	int sample(sample) ;
		sample:long_name = "Sample index" ;
		sample:units = "1" ;
		sample:comment = "Zero based index assigned to each sample period included in the file" ;
	int num_time_avg_ddms(num_time_avg_ddms) ;
		num_time_avg_ddms:long_name = "DDM index" ;
		num_time_avg_ddms:units = "1" ;
		num_time_avg_ddms:comment = "Additional dimension for those variables containing individual time-averaged values for each DDM contributing to the sample" ;
	byte ddm_source ;
		ddm_source:long_name = "DDM Source" ;
		ddm_source:units = "1" ;
		ddm_source:valid_range = 0b, 3b ;
		ddm_source:flag_values = 0b, 1b, 2b, 3b ;
		ddm_source:flag_meanings = "e2es gpss ddmi unknown" ;
		ddm_source:comment = "0=End-End Simulator (E2ES) 1=GPS signal simulator 2=CYGNSS DDMI 3=Source Unknown" ;
	byte spacecraft_num(sample) ;
		spacecraft_num:long_name = "Spacecraft Number" ;
		spacecraft_num:coordinates = "lat lon" ;
		spacecraft_num:units = "1" ;
		spacecraft_num:valid_min = 1 ;
		spacecraft_num:valid_max = 8 ;
		spacecraft_num:comment = "Numeric reference identifier (1-8) of the Cygnss spacecraft" ;
	byte spacecraft_id(sample) ;
		spacecraft_id:long_name = "Spacecraft Identifier" ;
		spacecraft_id:coordinates = "lat lon" ;
		spacecraft_id:units = "1" ;
		spacecraft_id:comment = "CCSDS Identifier (C-SCID) of the Cygnss spacecraft" ;
	byte prn_code(sample) ;
		prn_code:long_name = "GPS PRN code" ;
		prn_code:coordinates = "lat lon" ;
		prn_code:units = "1" ;
		prn_code:valid_min = 1 ;
		prn_code:valid_max = 32 ;
	byte antenna(sample) ;
		antenna:long_name = "Nadir Receive Antenna" ;
		antenna:coordinates = "lat lon" ;
		antenna:units = "1" ;
		antenna:valid_range = 2b, 3b ;
		antenna:flag_values = 2b, 3b ;
		antenna:flag_meanings = "nadir_starboard nadir_port" ;
		antenna:comment = "Nadir receive antenna associated with the retrieval" ;
	double sample_time(sample) ;
		sample_time:long_name = "Sample time " ;
		sample_time:standard_name = "time" ;
		sample_time:coordinates = "lat lon" ;
		sample_time:calendar = "gregorian" ;
		sample_time:comment = "Middle of the time averaging window, UTC" ;
		sample_time:units = "seconds since 2014-09-20 12:00:02.000000000" ;
	float lat(sample) ;
		lat:long_name = "latitude" ;
		lat:standard_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:comment = "Longitude of specular point of the DDM at the center of the time averaging window" ;
	float lon(sample) ;
		lon:long_name = "longitude" ;
		lon:standard_name = "longitude" ;
		lon:units = "degrees_east" ;
	float wind_speed(sample) ;
		wind_speed:long_name = "Wind Speed" ;
		wind_speed:standard_name = "wind_speed" ;
		wind_speed:coordinates = "lat lon" ;
		wind_speed:units = "m s-1" ;
		wind_speed:comment = "Time averaged retrieved wind speed" ;
	float wind_speed_error(sample) ;
		wind_speed_error:long_name = "Wind Speed Error" ;
		wind_speed_error:units = "m s-1" ;
		wind_speed_error:coordinates = "lat lon" ;
		wind_speed_error:comment = "Time averaged standard deviation of the error in retrieved wind speed" ;
	float mean_square_slope(sample) ;
		mean_square_slope:long_name = "Mean Square Slope" ;
		mean_square_slope:coordinates = "lat lon" ;
		mean_square_slope:units = "1" ;
		mean_square_slope:comment = "Time averaged mean square slope" ;
	float range_corr_gain(sample) ;
		range_corr_gain:long_name = "Range Corrected Gain" ;
		range_corr_gain:coordinates = "lat lon" ;
		range_corr_gain:units = "1e-27 meter-4" ;
		range_corr_gain:comment = "Time averaged RCG, calculated as RX-Antenna-gain/((R1^2)(R2^2))" ;
	float sig_wave_height(sample) ;
		sig_wave_height:long_name = "Significant Height of Wind and Swell Waves" ;
		sig_wave_height:standard_name = "sea_surface_wave_significant_height" ;
		sig_wave_height:coordinates = "lat lon" ;
		sig_wave_height:units = "meter" ;
		sig_wave_height:comment = "Significant wave height (SWH) at the location of the specular point of the DDM at the center of the time averaging window" ;
	float sea_surface_temp(sample) ;
		sea_surface_temp:long_name = "Sea Surface Temperature" ;
		sea_surface_temp:standard_name = "sea_surface_temperature" ;
		sea_surface_temp:coordinates = "lat lon" ;
		sea_surface_temp:units = "degree_Celsius" ;
		sea_surface_temp:comment = "SST at the location of the specular point of the DDM at the center of the time averaging window" ;
	float near_sea_surf_air_temp(sample) ;
		near_sea_surf_air_temp:long_name = "Near-surface Air Temperature (NAT)" ;
		near_sea_surf_air_temp:coordinates = "lat lon" ;
		near_sea_surf_air_temp:units = "degree_Celsius" ;
		near_sea_surf_air_temp:comment = "NAT at 2 meters at the location of the specular point of the DDM at the center of the time averaging window" ;
	float fresnel_reflec_coeff(sample) ;
		fresnel_reflec_coeff:long_name = "Fresnel reflection coefficient" ;
		fresnel_reflec_coeff:coordinates = "lat lon" ;
		fresnel_reflec_coeff:units = "1" ;
		fresnel_reflec_coeff:comment = "Fresnel reflection coefficient at the location of the specular point of the DDM at the center of the time averaging window" ;
	byte num_ddms(sample) ;
		num_ddms:long_name = "Number of DDMs" ;
		num_ddms:coordinates = "lat lon" ;
		num_ddms:units = "1" ;
		num_ddms:comment = "Actual number of DDMs that were time-averaged to produce wind retrieval" ;
	double ddm_time(sample, num_time_avg_ddms) ;
		ddm_time:long_name = "Level 1 DDM Times - UTC" ;
		ddm_time:standard_name = "time" ;
		ddm_time:coordinates = "ddm_lat ddm_lon" ;
		ddm_time:calendar = "gregorian" ;
		ddm_time:comment = "DDM timestamps (UTC) of each time-averaged DDM. Used together with the spacecraft Number and PRN code to look up Level 1 DDM Data" ;
		ddm_time:units = "seconds since 2014-09-20 12:00:02.000000000" ;
	float ddm_lat(sample, num_time_avg_ddms) ;
		ddm_lat:long_name = "DDM latitude" ;
		ddm_lat:standard_name = "latitude" ;
		ddm_lat:units = "degrees_north" ;
		ddm_lat:comment = "Location of specular point of each time-averaged DDM." ;
	float ddm_lon(sample, num_time_avg_ddms) ;
		ddm_lon:long_name = "DDM longitude" ;
		ddm_lon:standard_name = "longitude" ;
		ddm_lon:units = "degrees_east" ;
		ddm_lon:comment = "Location of specular point of each time-averaged DDM" ;
	float leading_edge_slope(sample, num_time_avg_ddms) ;
		leading_edge_slope:long_name = "DDM leading edge slope (LES) observable" ;
		leading_edge_slope:coordinates = "ddm_lat ddm_lon" ;
		leading_edge_slope:units = "1" ;
		leading_edge_slope:comment = "Leading edge slope for each time-averaged DDM." ;
	float ddm_area_avg(sample, num_time_avg_ddms) ;
		ddm_area_avg:long_name = "DDM area average (DDMA) observable" ;
		ddm_area_avg:coordinates = "ddm_lat ddm_lon" ;
		ddm_area_avg:units = "1" ;
		ddm_area_avg:comment = "DDM area for each time-averaged DDM." ;
	float wind_speed_from_les(sample, num_time_avg_ddms) ;
		wind_speed_from_les:long_name = "Wind speed derived from DDM LES" ;
		wind_speed_from_les:standard_name = "wind_speed" ;
		wind_speed_from_les:coordinates = "ddm_lat ddm_lon" ;
		wind_speed_from_les:units = "m s-1" ;
		wind_speed_from_les:comment = "Wind speed calculated from leading edge slope for each time-averaged DDM." ;
	float wind_speed_from_ddma(sample, num_time_avg_ddms) ;
		wind_speed_from_ddma:long_name = "Wind speed derived from DDM DDMA" ;
		wind_speed_from_ddma:standard_name = "wind_speed" ;
		wind_speed_from_ddma:coordinates = "ddm_lat ddm_lon" ;
		wind_speed_from_ddma:units = "m s-1" ;
		wind_speed_from_ddma:comment = "Wind speed calculated from DDM area for each time-averaged DDM." ;
	float ddm_wind_speed(sample, num_time_avg_ddms) ;
		ddm_wind_speed:long_name = "Wind speed - debiased and MV estimated" ;
		ddm_wind_speed:standard_name = "wind_speed" ;
		ddm_wind_speed:coordinates = "ddm_lat ddm_lon" ;
		ddm_wind_speed:units = "m s-1" ;
		ddm_wind_speed:comment = "Wind speed, debiased and MV-calculated, for each time-averaged DDM." ;
	float sp_incidence_angle(sample, num_time_avg_ddms) ;
		sp_incidence_angle:long_name = "Incidence angle of DDM specular point" ;
		sp_incidence_angle:coordinates = "ddm_lat ddm_lon" ;
		sp_incidence_angle:units = "degree" ;
		sp_incidence_angle:comment = "SP incidence angle for each time-averaged DDM, degrees from local vertical at location of specular point of DDM to line from specular point to CYGNSS spacecraft" ;
	float sp_azimuth_angle(sample, num_time_avg_ddms) ;
		sp_azimuth_angle:long_name = "Azimuth angle of DDM specular point" ;
		sp_azimuth_angle:coordinates = "ddm_lat ddm_lon" ;
		sp_azimuth_angle:units = "degree" ;
		sp_azimuth_angle:comment = "Azimuth angle of specular point for each time-averaged DDM, degrees from orbit frame +X axis to location of specular point of DDM" ;
	float ddm_range_corr_gain(sample) ;
		ddm_range_corr_gain:long_name = "Range Corrected Gains" ;
		ddm_range_corr_gain:coordinates = "lat lon" ;
		ddm_range_corr_gain:units = "1e-27 meter-4" ;
		ddm_range_corr_gain:comment = "RCG of each time-averaged DDM, calculated as RX-Antenna-gain-linear/((R1^2)(R2^2))" ;
	float sigma0(sample, num_time_avg_ddms) ;
		sigma0:long_name = "Sigma0" ;
		sigma0:coordinates = "ddm_lat ddm_lon" ;
		sigma0:units = "1" ;
		sigma0:comment = "BRCS normalized per scatter area for each time-averaged DDM" ;
	int sum_non_fatal_neg_wind_flags(sample) ;
		sum_non_fatal_neg_wind_flags:long_name = "Sum of non-fatal negative wind speed flags" ;
		sum_non_fatal_neg_wind_flags:coordinates = "lat lon" ;
		sum_non_fatal_neg_wind_flags:units = "1" ;
		sum_non_fatal_neg_wind_flags:comment = "DDM-level error flag, set if -5 <= DDM wind speed < 0 m/s" ;
	int sum_fatal_neg_wind_flags(sample) ;
		sum_fatal_neg_wind_flags:long_name = "Sum of fatal negative wind speed flags" ;
		sum_fatal_neg_wind_flags:coordinates = "lat lon" ;
		sum_fatal_neg_wind_flags:units = "1" ;
		sum_fatal_neg_wind_flags:comment = "DDM-level error flag, set if DDM wind speed < 5 m/s" ;
	int sum_non_fatal_high_wind_flags(sample) ;
		sum_non_fatal_high_wind_flags:long_name = "Sum of non-fatal high wind speed flags" ;
		sum_non_fatal_high_wind_flags:coordinates = "lat lon" ;
		sum_non_fatal_high_wind_flags:units = "1" ;
		sum_non_fatal_high_wind_flags:comment = "DDM-level error flag, set if 70 <= DDM wind speed < 100 m/s" ;
	int sum_fatal_high_wind_flags(sample) ;
		sum_fatal_high_wind_flags:long_name = "Sum of fatal high wind speed flags" ;
		sum_fatal_high_wind_flags:coordinates = "lat lon" ;
		sum_fatal_high_wind_flags:units = "1" ;
		sum_fatal_high_wind_flags:comment = "DDM-level error flag, set if DDM wind speed >= 100 m/s" ;
	int sum_neg_sigma0_ddma_area_flags(sample) ;
		sum_neg_sigma0_ddma_area_flags:long_name = "Sum of negative Sigma0 in DDMA area flags" ;
		sum_neg_sigma0_ddma_area_flags:coordinates = "lat lon" ;
		sum_neg_sigma0_ddma_area_flags:units = "1" ;
		sum_neg_sigma0_ddma_area_flags:comment = "DDM-level error flag, set if one or more Sigma0 DDM bins in the DDMA area are negative" ;
	int sum_low_range_corr_gain_flags(sample) ;
		sum_low_range_corr_gain_flags:long_name = "Sum of low Range Corrected gain flags" ;
		sum_low_range_corr_gain_flags:coordinates = "lat lon" ;
		sum_low_range_corr_gain_flags:units = "1" ;
		sum_low_range_corr_gain_flags:comment = "DDM-level error flag, set if DDM range corrected gain < 3" ;
	int sum_high_sp_incidence_angle_flags(sample) ;
		sum_high_sp_incidence_angle_flags:long_name = "Sum of high specular point incidence angle flags" ;
		sum_high_sp_incidence_angle_flags:coordinates = "lat lon" ;
		sum_high_sp_incidence_angle_flags:units = "1" ;
		sum_high_sp_incidence_angle_flags:comment = "DDM-Level error flag, set if DDM specular point incidence angle > 70" ;
	int sum_ddma_area_near_edge_flags(sample) ;
		sum_ddma_area_near_edge_flags:long_name = "Sum of DDMA area near edge of DDM flags" ;
		sum_ddma_area_near_edge_flags:coordinates = "lat lon" ;
		sum_ddma_area_near_edge_flags:units = "1" ;
		sum_ddma_area_near_edge_flags:comment = "DDM-level error flag, set if any edge of the DDMA area coincides with an edge of the DDM" ;
	int sum_sp_outside_ddma_area_flags(sample) ;
		sum_sp_outside_ddma_area_flags:long_name = "Sum of specular point outside the edge of DDMA area flags" ;
		sum_sp_outside_ddma_area_flags:coordinates = "lat lon" ;
		sum_sp_outside_ddma_area_flags:units = "1" ;
		sum_sp_outside_ddma_area_flags:comment = "DDM-level error flag, set if any part of the DDMA area falls outside of the DDM" ;
	int sum_l1_poor_overall_quality_flags(sample) ;
		sum_l1_poor_overall_quality_flags:long_name = "Sum of L1 DDM poor overall quality flags" ;
		sum_l1_poor_overall_quality_flags:coordinates = "lat lon" ;
		sum_l1_poor_overall_quality_flags:units = "1" ;
		sum_l1_poor_overall_quality_flags:comment = "This flag is copied directly from the L1 input file. It indicates that L1 processing determined that the DDM was of poor overall quality." ;

// global attributes:
		:Conventions = "CF-1.6, ACDD-1.3, ISO-8601" ;
		:standard_name_vocabulary = "CF Standard Name Table v30" ;
		:project = "CYGNSS" ;
		:summary = "TBD. Per ACDD, a paragraph analogous to an abstract." ;
		:processing_level = "Time-tagged, precision geolocated average windspeed and mean square slope of 25x25Km cells centered on specular points and associated metadata." ;
		:comment = "L1 DDMs are processed to produce windspeed and mean square slope" ;
		:creator_type = "institution" ;
		:institution = "University of Michigan Space Physics Research Lab (SPRL)" ;
		:creator_name = "CYGNSS Science Operations Center" ;
		:publisher_name = "PO.DAAC" ;
		:publisher_email = "podaac@podaac.jpl.nasa.gov" ;
		:publisher_url = "​http://podaac.jpl.nasa.gov" ;
		:sensor = "Delay Doppler Mapping Instrument (DDMI)" ;
		:source = "Delay Doppler maps (DDM) obtained from the DDMI aboard CYGNSS observatory constellation" ;
		:program = "TBD. Per ACDD: <<<The overarching program(s) of which the dataset is a part. A program consists of a set (or portfolio) of related and possibly interdependent projects that meet an overarching objective. Examples: \'GHRSST\', \'NOAA CDR\', \'NASA EOS\', \'JPSS\', \'GOES-R\'.>>>" ;
		:references = "TBD. Per ACDD: <<<Published or web-based references that describe the data or methods used to produce it. Recommend URIs (such as a URL or DOI) for papers or other references.>>>" ;
		:version_id = "1.0" ;
		:title = "CYGNSS Level 2 Science Data Record Version 1.0" ;
		:ShortName = "CYGNSS_L2_V1.0" ;
		:id = "PODAAC-CYGNS-L2X10" ;
		:netcdf_version_id = "4.3.3.1 of Dec 10 2015 16:44:18 $" ;
		:date_created = "2016-06-16T13:04:54Z" ;
		:date_issued = "2016-06-16T13:04:54Z" ;
		:history = "Thu Jun 16 13:05:00 2016: ncks -O -L1 -a /tmp/qt_temp.T16106 out.nc\n./produce-L2-files /home/butlerti/data/l0_csv_tests/June9_2016_a.nc --output-file out.nc" ;
		:time_coverage_resolution = "P0DT0H0M1S" ;
		:time_coverage_start = "2014-09-20T12:00:02.000000000Z" ;
		:time_coverage_end = "2014-09-20T13:40:00.000000000Z" ;
		:time_coverage_duration = "P0DT1H39M59S" ;
		:l2_algorithm_version = "1" ;
		:ddma_les_sel_lookup_tables_version = "2" ;
		:time_averaging_lookup_tables_version = "1" ;
		:ddma_wind_lookup_tables_version = "5" ;
		:les_wind_lookup_tables_version = "5" ;
		:covariance_lookup_tables_version = "2" ;
		:standard_deviation_lookup_tables_version = "2" ;
		:geospatial_lat_min = "-54.606N" ;
		:geospatial_lat_max = "51.601N" ;
		:geospatial_lon_min = "40.094E" ;
		:geospatial_lon_max = "355.607E" ;
		:NCO = "4.4.4" ;
}
