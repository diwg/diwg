netcdf S5P_OFFL_L2__AER_AI_20070813T033313_20070813T051437_04226_01_000900_20151102T000000 {

// global attributes:
		:time_reference = "2007-08-13T00:00:00Z" ;
		:time_reference_days_since_1950 = 21043 ;
		:time_reference_julian_day = 2454325.5 ;
		:time_reference_seconds_since_1970 = 1186963200L ;
		:time_coverage_start = "2007-08-13T03:33:13Z" ;
		:time_coverage_end = "2007-08-13T05:14:37Z" ;
		:time_coverage_duration = "PT6084.000S" ;
		:time_coverage_resolution = "PT10.294S" ;

group: PRODUCT {
  dimensions:
  	scanline = UNLIMITED ; // (592 currently)
  	ground_pixel = 316 ;
  	corner = 4 ;
  	time = 1 ;
  variables:
  	int scanline(scanline) ;
  		scanline:units = "1" ;
  		scanline:long_name = "along-track dimension index" ;
  		scanline:comment = "This coordinate variable defines the indices along track; index starts at 0" ;
  		scanline:_FillValue = -2147483647 ;
  	int ground_pixel(ground_pixel) ;
  		ground_pixel:units = "1" ;
  		ground_pixel:long_name = "across-track dimension index" ;
  		ground_pixel:comment = "This coordinate variable defines the indices across track, from west to east; index starts at 0" ;
  		ground_pixel:_FillValue = -2147483647 ;
  	int time(time) ;
  		time:units = "seconds since 2010-01-01 00:00:00" ;
  		time:standard_name = "time" ;
  		time:long_name = "reference time for the measurements" ;
  		time:comment = "The time in this variable corresponds to the time in the time_reference global attribute" ;
  		time:_FillValue = -2147483647 ;
  	int corner(corner) ;
  		corner:units = "1" ;
  		corner:long_name = "pixel corner index" ;
  		corner:comment = "This coordinate variable defines the indices for the pixel corners; index starts at 0 (counter-clockwise, starting from south-western corner of the pixel in ascending part of the orbit)" ;
  		corner:_FillValue = -2147483647 ;
  	float latitude(time, scanline, ground_pixel) ;
  		latitude:long_name = "pixel center latitude" ;
  		latitude:units = "degrees_north" ;
  		latitude:standard_name = "latitude" ;
  		latitude:valid_min = -90.f ;
  		latitude:valid_max = 90.f ;
  		latitude:bounds = "/PRODUCT/SUPPORT_DATA/GEOLOCATIONS/latitude_bounds" ;
  		latitude:_FillValue = 9.96921e+36f ;
  	float longitude(time, scanline, ground_pixel) ;
  		longitude:long_name = "pixel center longitude" ;
  		longitude:units = "degrees_east" ;
  		longitude:standard_name = "longitude" ;
  		longitude:valid_min = -180.f ;
  		longitude:valid_max = 180.f ;
  		longitude:bounds = "/PRODUCT/SUPPORT_DATA/GEOLOCATIONS/longitude_bounds" ;
  		longitude:_FillValue = 9.96921e+36f ;
  	int delta_time(time, scanline) ;
  		delta_time:long_name = "offset from reference start time of measurement" ;
  		delta_time:units = "milliseconds" ;
  		delta_time:_FillValue = -2147483647 ;
  	string time_utc(time, scanline) ;
  		time_utc:long_name = "Time of observation as ISO 8601 date-time string" ;
  		string time_utc:_FillValue = "" ;
  	float aerosol_index_354_388(time, scanline, ground_pixel) ;
  		aerosol_index_354_388:units = "1" ;
  		aerosol_index_354_388:standard_name = "ultraviolet_aerosol_index" ;
  		aerosol_index_354_388:comment = "Aerosol index from 388 and 354 nm" ;
  		aerosol_index_354_388:long_name = "Aerosol index from 388 and 354 nm" ;
  		aerosol_index_354_388:radiation_wavelength = 354.f, 388.f ;
  		aerosol_index_354_388:coordinates = "longitude latitude" ;
  		aerosol_index_354_388:ancillary_variables = "aerosol_index_354_388_precision" ;
  		aerosol_index_354_388:_FillValue = 9.96921e+36f ;
  	float aerosol_index_354_388_precision(time, scanline, ground_pixel) ;
  		aerosol_index_354_388_precision:units = "1" ;
  		aerosol_index_354_388_precision:standard_name = "ultraviolet_aerosol_index standard_error" ;
  		aerosol_index_354_388_precision:comment = "Precision of aerosol index from 388 and 354 nm" ;
  		aerosol_index_354_388_precision:long_name = "Precision of aerosol index from 388 and 354 nm" ;
  		aerosol_index_354_388_precision:radiation_wavelength = 354.f, 388.f ;
  		aerosol_index_354_388_precision:coordinates = "longitude latitude" ;
  		aerosol_index_354_388_precision:_FillValue = 9.96921e+36f ;

  group: SUPPORT_DATA {

    group: GEOLOCATIONS {
      variables:
      	float satellite_latitude(time, scanline) ;
      		satellite_latitude:long_name = "sub satellite latitude" ;
      		satellite_latitude:units = "degrees_north" ;
      		satellite_latitude:comment = "Latitude of the geodetic sub satellite point on the WGS84 reference ellipsoid" ;
      		satellite_latitude:valid_min = -90.f ;
      		satellite_latitude:valid_max = 90.f ;
      		satellite_latitude:_FillValue = 9.96921e+36f ;
      	float satellite_longitude(time, scanline) ;
      		satellite_longitude:long_name = "satellite_longitude" ;
      		satellite_longitude:units = "degrees_east" ;
      		satellite_longitude:comment = "Longitude of the geodetic sub satellite point on the WGS84 reference ellipsoid" ;
      		satellite_longitude:valid_min = -180.f ;
      		satellite_longitude:valid_max = 180.f ;
      		satellite_longitude:_FillValue = 9.96921e+36f ;
      	float satellite_altitude(time, scanline) ;
      		satellite_altitude:long_name = "satellite altitude" ;
      		satellite_altitude:units = "m" ;
      		satellite_altitude:comment = "The altitude of the satellite with respect to the geodetic sub satellite point on the WGS84 reference ellipsoid" ;
      		satellite_altitude:valid_min = 700000.f ;
      		satellite_altitude:valid_max = 900000.f ;
      		satellite_altitude:_FillValue = 9.96921e+36f ;
      	float satellite_orbit_phase(time, scanline) ;
      		satellite_orbit_phase:long_name = "fractional satellite orbit phase" ;
      		satellite_orbit_phase:units = "1" ;
      		satellite_orbit_phase:comment = "Relative offset [0.0, ..., 1.0] of the measurement in the orbit" ;
      		satellite_orbit_phase:valid_min = -0.02f ;
      		satellite_orbit_phase:valid_max = 1.02f ;
      		satellite_orbit_phase:_FillValue = 9.96921e+36f ;
      	float solar_zenith_angle(time, scanline, ground_pixel) ;
      		solar_zenith_angle:long_name = "solar zenith angle" ;
      		solar_zenith_angle:standard_name = "solar_zenith_angle" ;
      		solar_zenith_angle:units = "degree" ;
      		solar_zenith_angle:valid_min = 0.f ;
      		solar_zenith_angle:valid_max = 180.f ;
      		solar_zenith_angle:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		solar_zenith_angle:comment = "Solar zenith angle at the ground pixel location on the reference ellipsoid. Angle is measured away from the vertical" ;
      		solar_zenith_angle:_FillValue = 9.96921e+36f ;
      	float solar_azimuth_angle(time, scanline, ground_pixel) ;
      		solar_azimuth_angle:long_name = "solar azimuth angle" ;
      		solar_azimuth_angle:standard_name = "solar_azimuth_angle" ;
      		solar_azimuth_angle:units = "degree" ;
      		solar_azimuth_angle:valid_min = 0.f ;
      		solar_azimuth_angle:valid_max = 360.f ;
      		solar_azimuth_angle:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		solar_azimuth_angle:comment = "Solar azimuth angle at the ground pixel location on the reference ellipsoid. Angle is measured clockwise from the North (East = 90, South = 180, West = 270)" ;
      		solar_azimuth_angle:_FillValue = 9.96921e+36f ;
      	float viewing_zenith_angle(time, scanline, ground_pixel) ;
      		viewing_zenith_angle:long_name = "viewing zenith angle" ;
      		viewing_zenith_angle:standard_name = "viewing_zenith_angle" ;
      		viewing_zenith_angle:units = "degree" ;
      		viewing_zenith_angle:valid_min = 0.f ;
      		viewing_zenith_angle:valid_max = 180.f ;
      		viewing_zenith_angle:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		viewing_zenith_angle:comment = "Zenith angle of the satellite at the ground pixel location on the reference ellipsoid. Angle is measured away from the vertical" ;
      		viewing_zenith_angle:_FillValue = 9.96921e+36f ;
      	float viewing_azimuth_angle(time, scanline, ground_pixel) ;
      		viewing_azimuth_angle:long_name = "viewing azimuth angle" ;
      		viewing_azimuth_angle:standard_name = "viewing_azimuth_angle" ;
      		viewing_azimuth_angle:units = "degree" ;
      		viewing_azimuth_angle:valid_min = 0.f ;
      		viewing_azimuth_angle:valid_max = 360.f ;
      		viewing_azimuth_angle:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		viewing_azimuth_angle:comment = "Satellite azimuth angle at the ground pixel location on the reference ellipsoid. Angle is measured clockwise from the North (East = 90, South = 180, West = 270)" ;
      		viewing_azimuth_angle:_FillValue = 9.96921e+36f ;
      	float latitude_bounds(time, scanline, ground_pixel, corner) ;
      		latitude_bounds:_FillValue = 9.96921e+36f ;
      	float longitude_bounds(time, scanline, ground_pixel, corner) ;
      		longitude_bounds:_FillValue = 9.96921e+36f ;
      } // group GEOLOCATIONS

    group: DETAILED_RESULTS {
      variables:
      	uint processing_quality_flags(time, scanline, ground_pixel) ;
      		processing_quality_flags:long_name = "Processing quality flags" ;
      		processing_quality_flags:comment = "Flags indicating conditions that affect quality of the retrieval." ;
      		processing_quality_flags:flag_meanings = "success radiance_missing irradiance_missing input_spectrum_missing reflectance_range_error ler_range_error snr_range_error sza_range_error vza_range_error lut_range_error ozone_range_error wavelength_offset_error initialization_error memory_error assertion_error io_error numerical_error lut_error ISRF_error convergence_error cloud_filter_convergence_error max_iteration_convergence_error aot_lower_boundary_convergence_error other_boundary_convergence_error geolocation_error ch4_noscat_zero_error h2o_noscat_zero_error max_optical_thickness_error aerosol_boundary_error boundary_hit_error chi2_error svd_error dfs_error radiative_transfer_error optimal_estimation_error profile_error cloud_error model_error number_of_input_data_points_too_low_error cloud_pressure_spread_too_low_error cloud_too_low_level_error generic_range_error generic_exception input_spectrum_alignment_error abort_error wrong_input_type_error wavelength_calibration_error coregistration_error solar_eclipse_filter cloud_filter altitude_consistency_filter altitude_roughness_filter sun_glint_filter mixed_surface_type_filter snow_ice_filter aai_filter cloud_fraction_fresco_filter aai_scene_albedo_filter small_pixel_radiance_std_filter cloud_fraction_viirs_filter cirrus_reflectance_viirs_filter cf_viirs_swir_ifov_filter cf_viirs_swir_ofova_filter cf_viirs_swir_ofovb_filter cf_viirs_swir_ofovc_filter cf_viirs_nir_ifov_filter cf_viirs_nir_ofova_filter cf_viirs_nir_ofovb_filter cf_viirs_nir_ofovc_filter refl_cirrus_viirs_swir_filter refl_cirrus_viirs_nir_filter diff_refl_cirrus_viirs_filter ch4_noscat_ratio_filter ch4_noscat_ratio_std_filter h2o_noscat_ratio_filter h2o_noscat_ratio_std_filter diff_psurf_fresco_ecmwf_filter psurf_fresco_stdv_filter ocean_filter time_range_filter pixel_or_scanline_index_filter geographic_region_filter input_spectrum_warning wavelength_calibration_warning extrapolation_warning sun_glint_warning south_atlantic_anomaly_warning sun_glint_correction snow_ice_warning cloud_warning AAI_warning pixel_level_input_data_missing data_range_warning low_cloud_fraction_warning altitude_consistency_warning signal_to_noise_ratio_warning deconvolution_warning so2_volcanic_origin_likely_warning so2_volcanic_origin_certain_warning interpolation_warning" ;
      		processing_quality_flags:flag_masks = 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 256U, 512U, 1024U, 2048U, 4096U, 8192U, 16384U, 32768U, 65536U, 131072U, 262144U, 524288U, 1048576U, 2097152U, 4194304U, 8388608U, 16777216U, 33554432U ;
      		processing_quality_flags:flag_values = 0U, 1U, 2U, 3U, 4U, 5U, 6U, 7U, 8U, 9U, 10U, 11U, 12U, 13U, 14U, 15U, 16U, 17U, 18U, 19U, 20U, 21U, 22U, 23U, 24U, 25U, 26U, 27U, 28U, 29U, 30U, 31U, 32U, 33U, 34U, 35U, 36U, 37U, 38U, 39U, 40U, 41U, 42U, 43U, 44U, 45U, 46U, 47U, 64U, 65U, 66U, 67U, 68U, 69U, 70U, 71U, 72U, 73U, 74U, 75U, 76U, 77U, 78U, 79U, 80U, 81U, 82U, 83U, 84U, 85U, 86U, 87U, 88U, 89U, 90U, 91U, 92U, 93U, 94U, 95U, 96U, 97U, 256U, 512U, 1024U, 2048U, 4096U, 8192U, 16384U, 32768U, 65536U, 131072U, 262144U, 524288U, 1048576U, 2097152U, 4194304U, 8388608U, 16777216U, 33554432U ;
      		processing_quality_flags:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		processing_quality_flags:_FillValue = 4294967295U ;
      	ushort number_of_spectral_points_in_retrieval(time, scanline, ground_pixel) ;
      		number_of_spectral_points_in_retrieval:long_name = "number of spectral points used in the retrieval." ;
      		number_of_spectral_points_in_retrieval:comment = "Flags indicating conditions that affect quality of the retrieval." ;
      		number_of_spectral_points_in_retrieval:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		number_of_spectral_points_in_retrieval:_FillValue = 65535US ;
      	float scene_albedo_388(time, scanline, ground_pixel) ;
      		scene_albedo_388:units = "1" ;
      		scene_albedo_388:long_name = "Scene albedo at 388 nm calculated from the top of atmosphere reflectance. For a cloud- and aerosol-free scene this is equivalent to the surface albedo" ;
      		scene_albedo_388:radiation_wavelength = 388.f ;
      		scene_albedo_388:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		scene_albedo_388:ancillary_variables = "scene_albedo_388_precision" ;
      		scene_albedo_388:_FillValue = 9.96921e+36f ;
      	float scene_albedo_388_precision(time, scanline, ground_pixel) ;
      		scene_albedo_388_precision:units = "1" ;
      		scene_albedo_388_precision:long_name = "Precision of the scene albedo at 388 nm calculated from the top of atmosphere reflectance and its precision. For a cloud- and aerosol-free scene this is equivalent to the surface albedo" ;
      		scene_albedo_388_precision:radiation_wavelength = 388.f ;
      		scene_albedo_388_precision:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		scene_albedo_388_precision:_FillValue = 9.96921e+36f ;
      	float reflectance_measured_354(time, scanline, ground_pixel) ;
      		reflectance_measured_354:units = "1" ;
      		reflectance_measured_354:standard_name = "toa_bidirectional_reflectance" ;
      		reflectance_measured_354:long_name = "Top of atmosphere reflectance at 354 nm" ;
      		reflectance_measured_354:radiation_wavelength = 354.f ;
      		reflectance_measured_354:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		reflectance_measured_354:ancillary_variables = "reflectance_measured_354_precision" ;
      		reflectance_measured_354:_FillValue = 9.96921e+36f ;
      	float reflectance_measured_354_precision(time, scanline, ground_pixel) ;
      		reflectance_measured_354_precision:units = "1" ;
      		reflectance_measured_354_precision:standard_name = "toa_bidirectional_reflectance standard_error" ;
      		reflectance_measured_354_precision:long_name = "Precision of the top of atmosphere reflectance at 354 nm" ;
      		reflectance_measured_354_precision:radiation_wavelength = 354.f ;
      		reflectance_measured_354_precision:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		reflectance_measured_354_precision:_FillValue = 9.96921e+36f ;
      	float reflectance_measured_388(time, scanline, ground_pixel) ;
      		reflectance_measured_388:units = "1" ;
      		reflectance_measured_388:standard_name = "toa_bidirectional_reflectance" ;
      		reflectance_measured_388:long_name = "Top of atmosphere reflectance at 388 nm" ;
      		reflectance_measured_388:radiation_wavelength = 388.f ;
      		reflectance_measured_388:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		reflectance_measured_388:ancillary_variables = "reflectance_measured_388_precision" ;
      		reflectance_measured_388:_FillValue = 9.96921e+36f ;
      	float reflectance_measured_388_precision(time, scanline, ground_pixel) ;
      		reflectance_measured_388_precision:units = "1" ;
      		reflectance_measured_388_precision:standard_name = "toa_bidirectional_reflectance standard_error" ;
      		reflectance_measured_388_precision:long_name = "Precision of the top of atmosphere reflectance at 388 nm" ;
      		reflectance_measured_388_precision:radiation_wavelength = 388.f ;
      		reflectance_measured_388_precision:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		reflectance_measured_388_precision:_FillValue = 9.96921e+36f ;
      	float reflectance_calculated_354(time, scanline, ground_pixel) ;
      		reflectance_calculated_354:units = "1" ;
      		reflectance_calculated_354:standard_name = "toa_bidirectional_reflectance" ;
      		reflectance_calculated_354:long_name = "Calculated top of atmosphere reflectance at 354 nm" ;
      		reflectance_calculated_354:radiation_wavelength = 354.f ;
      		reflectance_calculated_354:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		reflectance_calculated_354:ancillary_variables = "reflectance_calculated_354_precision" ;
      		reflectance_calculated_354:_FillValue = 9.96921e+36f ;
      	float reflectance_calculated_354_precision(time, scanline, ground_pixel) ;
      		reflectance_calculated_354_precision:units = "1" ;
      		reflectance_calculated_354_precision:standard_name = "toa_bidirectional_reflectance standard_error" ;
      		reflectance_calculated_354_precision:long_name = "Precision of the calculated top of atmosphere reflectance at 354 nm" ;
      		reflectance_calculated_354_precision:radiation_wavelength = 354.f ;
      		reflectance_calculated_354_precision:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		reflectance_calculated_354_precision:_FillValue = 9.96921e+36f ;
      	float wavelength_calibration_offset(time, scanline, ground_pixel) ;
      		wavelength_calibration_offset:long_name = "wavelength offset" ;
      		wavelength_calibration_offset:units = "nm" ;
      		wavelength_calibration_offset:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		wavelength_calibration_offset:ancillary_variables = "wavelength_calibration_offset_precision" ;
      		wavelength_calibration_offset:comment = "true wavelength = nominal wavelength + wavelength offset + wavelength stretch * scaled wavelength" ;
      		wavelength_calibration_offset:_FillValue = 9.96921e+36f ;
      		wavelength_calibration_offset:wavelength_fit_window_start = 338. ;
      		wavelength_calibration_offset:wavelength_fit_window_end = 390. ;
      	float wavelength_calibration_offset_precision(time, scanline, ground_pixel) ;
      		wavelength_calibration_offset_precision:long_name = "wavelength offset precision" ;
      		wavelength_calibration_offset_precision:units = "nm" ;
      		wavelength_calibration_offset_precision:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		wavelength_calibration_offset_precision:_FillValue = 9.96921e+36f ;
      	float wavelength_calibration_chi_squared(time, scanline, ground_pixel) ;
      		wavelength_calibration_chi_squared:long_name = "wavelength calibration chi squared" ;
      		wavelength_calibration_chi_squared:units = "1" ;
      		wavelength_calibration_chi_squared:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		wavelength_calibration_chi_squared:_FillValue = 9.96921e+36f ;
      } // group DETAILED_RESULTS

    group: INPUT_DATA {
      variables:
      	float surface_altitude(time, scanline, ground_pixel) ;
      		surface_altitude:long_name = "surface altitude" ;
      		surface_altitude:standard_name = "surface_altitude" ;
      		surface_altitude:units = "m" ;
      		surface_altitude:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		surface_altitude:source = "http://topotools.cr.usgs.gov/gmted_viewer/" ;
      		surface_altitude:comment = "The mean of the sub-pixels of the surface altitude above the reference geoid (WGS84) within the approximate field of view, based on the GMTED2010 surface elevation database" ;
      		surface_altitude:_FillValue = 9.96921e+36f ;
      	float surface_altitude_precision(time, scanline, ground_pixel) ;
      		surface_altitude_precision:long_name = "surface altitude precision" ;
      		surface_altitude_precision:standard_name = "surface_altitude standard_error" ;
      		surface_altitude_precision:units = "m" ;
      		surface_altitude_precision:standard_error_multiplier = 1.f ;
      		surface_altitude_precision:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		surface_altitude_precision:source = "http://topotools.cr.usgs.gov/gmted_viewer/" ;
      		surface_altitude_precision:comment = "The standard deviation of sub-pixels used in calculating the mean surface altitude above the reference geoid (WGS84) within the approximate field of view, based on the GMTED2010 surface elevation database" ;
      		surface_altitude_precision:_FillValue = 9.96921e+36f ;
      	ubyte surface_classification(time, scanline, ground_pixel) ;
      		surface_classification:long_name = "land-water mask" ;
      		surface_classification:comment = "flag indicating land/water and further surface classifications for the ground pixel" ;
      		surface_classification:source = "USGS (http://edc2.usgs.gov/glcc/globdoc2_0.php) and NASA SDP toolkit (http://newsroom.gsfc.nasa.gov/sdptoolkit/toolkit.html)" ;
      		surface_classification:flag_meanings = "land, water, some_water, coast, value_covers_majority_of_pixel, water+shallow_ocean, water+shallow_inland_water, water+ocean_coastline-lake_shoreline, water+intermittent_water, water+deep_inland_water, water+continental_shelf_ocean, water+deep_ocean, land+urban_and_built-up_land, land+dryland_cropland_and_pasture, land+irrigated_cropland_and_pasture, land+mixed_dryland-irrigated_cropland_and_pasture, land+cropland-grassland_mosaic, land+cropland-woodland_mosaic, land+grassland, land+shrubland, land+mixed_shrubland-grassland, land+savanna, land+deciduous_broadleaf_forest, land+deciduous_needleleaf_forest, land+evergreen_broadleaf_forest, land+evergreen_needleleaf_forest, land+mixed_forest, land+herbaceous_wetland, land+wooded_wetland, land+barren_or_sparsely_vegetated, land+herbaceous_tundra, land+wooded_tundra, land+mixed_tundra, land+bare_ground_tundra, land+snow_or_ice" ;
      		surface_classification:flag_values = 0UB, 1UB, 2UB, 3UB, 4UB, 9UB, 17UB, 25UB, 33UB, 41UB, 49UB, 57UB, 8UB, 16UB, 24UB, 32UB, 40UB, 48UB, 56UB, 64UB, 72UB, 80UB, 88UB, 96UB, 104UB, 112UB, 120UB, 128UB, 136UB, 144UB, 152UB, 160UB, 168UB, 176UB, 184UB ;
      		surface_classification:flag_masks = 3UB, 3UB, 3UB, 3UB, 4UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB ;
      		surface_classification:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		surface_classification:_FillValue = 255UB ;
      	float small_pixel_variance(time, scanline, ground_pixel) ;
      		small_pixel_variance:long_name = "scaled small pixel variance" ;
      		small_pixel_variance:units = "1" ;
      		small_pixel_variance:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		small_pixel_variance:comment = "The variance of the reflectances of the small pixels" ;
      		small_pixel_variance:_FillValue = 9.96921e+36f ;
      		small_pixel_variance:radiation_wavelength = 9.96921e+36f ;
      	float O3_total_vertical_column(time, scanline, ground_pixel) ;
      		O3_total_vertical_column:units = "mol m-2" ;
      		O3_total_vertical_column:standard_name = "atmosphere_mole_content_of_ozone" ;
      		O3_total_vertical_column:long_name = "total column amount of ozone" ;
      		O3_total_vertical_column:source = "" ;
      		O3_total_vertical_column:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		O3_total_vertical_column:multiplication_factor_to_convert_to_DU = 2241.15f ;
      		O3_total_vertical_column:multiplication_factor_to_convert_to_molecules_percm2 = 6.022141e+19f ;
      		O3_total_vertical_column:_FillValue = 9.96921e+36f ;
      	float surface_pressure(time, scanline, ground_pixel) ;
      		surface_pressure:units = "hPa" ;
      		surface_pressure:standard_name = "surface_air_pressure" ;
      		surface_pressure:long_name = "surface_air_pressure" ;
      		surface_pressure:source = "" ;
      		surface_pressure:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		surface_pressure:_FillValue = 9.96921e+36f ;
      } // group INPUT_DATA
    } // group SUPPORT_DATA
  } // group PRODUCT

group: METADATA {

  group: QA_STATISTICS {
    dimensions:
    	vertices = 2 ;
    	aerosol_index_354_388_histogram_axis = 100 ;
    	aerosol_index_354_388_pdf_axis = 400 ;
    	aerosol_index_340_380_histogram_axis = 100 ;
    	aerosol_index_340_380_pdf_axis = 400 ;
    variables:
    	float aerosol_index_354_388_histogram_axis(aerosol_index_354_388_histogram_axis) ;
    		aerosol_index_354_388_histogram_axis:units = "1" ;
    		aerosol_index_354_388_histogram_axis:comment = "Histogram axis of the aerosol index" ;
    		aerosol_index_354_388_histogram_axis:long_name = "Histogram axis of the aerosol index" ;
    		aerosol_index_354_388_histogram_axis:bounds = "aerosol_index_354_388_histogram_bounds" ;
    		aerosol_index_354_388_histogram_axis:_FillValue = 9.96921e+36f ;
    	float aerosol_index_354_388_histogram_bounds(aerosol_index_354_388_histogram_axis, vertices) ;
    		aerosol_index_354_388_histogram_bounds:_FillValue = 9.96921e+36f ;
    	int aerosol_index_354_388_histogram(aerosol_index_340_380_histogram_axis) ;
    		aerosol_index_354_388_histogram:comment = "Histogram of the aerosol index of the 354/388 nm pair in the current granule" ;
    		aerosol_index_354_388_histogram:_FillValue = -2147483647 ;
    		aerosol_index_354_388_histogram:number_of_overflow_values = 0 ;
    		aerosol_index_354_388_histogram:number_of_underflow_values = 3 ;

    // group attributes:
    		:number_of_groundpixels = 187072 ;
    		:number_of_processed_pixels = 14208 ;
    		:number_of_successfully_processed_pixels = 11348 ;
    		:number_of_rejected_pixels_not_enough_spectrum = 0 ;
    		:number_of_failed_retrievals = 2860 ;
    		:number_of_ground_pixels_with_warnings = 761 ;
    } // group QA_STATISTICS

  group: ALGORITHM_SETTINGS {

    // group attributes:
    		:algo.algorithm_variant = "1" ;
    		:algo.n_pair = "2" ;
    		:algo.pair_1.delta_wavelength = "1" ;
    		:algo.pair_1.id = "OMI_pair" ;
    		:algo.pair_1.min_wavelength = "1" ;
    		:algo.pair_1.number_spectral_pixels = "5" ;
    		:algo.pair_1.wavelength_1 = "354" ;
    		:algo.pair_1.wavelength_2 = "388" ;
    		:input.1.band = "3" ;
    		:input.1.irrType = "L1B_IR_UVN" ;
    		:input.1.type = "L1B_RA_BD3" ;
    		:input.count = "1" ;
    		:output.1.band = "3" ;
    		:output.1.config = "cfg/product/product.AER_AI.xml" ;
    		:output.1.type = "L2__AER_AI" ;
    		:output.count = "1" ;
    		:output.histogram.aerosol_index_354_388.end = "14" ;
    		:output.histogram.aerosol_index_354_388.start = "-6" ;
    		:processing.algorithm = "AER_AI" ;
    		:processing.szaMax = "88.0" ;
    		:wavelength_calibration.convergance_threshold = "1." ;
    		:wavelength_calibration.include_ring = "yes" ;
    		:wavelength_calibration.initial_guess.a0 = "1.0" ;
    		:wavelength_calibration.initial_guess.a1 = "0.1" ;
    		:wavelength_calibration.initial_guess.a2 = "0.01" ;
    		:wavelength_calibration.initial_guess.ring = "0.06" ;
    		:wavelength_calibration.initial_guess.shift = "0.0" ;
    		:wavelength_calibration.max_iterations = "12" ;
    		:wavelength_calibration.perform_wavelength_fit = "yes" ;
    		:wavelength_calibration.polynomial_order = "3" ;
    		:wavelength_calibration.sigma.a0 = "1.0" ;
    		:wavelength_calibration.sigma.a1 = "0.1" ;
    		:wavelength_calibration.sigma.ring = "0.06" ;
    		:wavelength_calibration.window = "338.0, 390.0" ;
    } // group ALGORITHM_SETTINGS

  group: GRANULE_DESCRIPTION {

    // group attributes:
    		:InstrumentName = "TROPOMI" ;
    		:MissionName = "Sentinel-5 precursor" ;
    		:MissionShortName = "S5P" ;
    		:ProcessLevel = "2" ;
    		:ProductFormatVersion = 1 ;
    		:ProductShortName = "L2__AER_AI" ;
    		:GranuleStart = "2007-08-13T03:33:13Z" ;
    		:GranuleEnd = "2007-08-13T05:14:37Z" ;
    		:ProcessingCenter = "KNMI" ;
    		:ProcessingNode = "bhltrdl2.knmi.nl" ;
    		:ProcessorVersion = "0.9.0" ;
    		:ProcessingMode = "Offline" ;
    } // group GRANULE_DESCRIPTION

  group: ESA_METADATA {

    group: earth_explorer_header {

      // group attributes:
      		:objectType = "Earth_Explorer_Header" ;

      group: fixed_header {

        // group attributes:
        		:objectType = "Fixed_Header" ;
        		:Notes = "" ;
        		:Mission = "S5P" ;
        		:File_Name = "S5P_OFFL_L2__AER_AI_20070813T033313_20070813T051437_04226_01_000900_20151102T000000" ;
        		:File_Description = "Aerosol index with a spatial resolution of 7x7km2 observed at about 13:30 local solar time from spectra measured by TROPOMI" ;
        		:File_Class = "OFFL" ;
        		:File_Type = "L2__AER_AI" ;
        		:File_Version = 1 ;

        group: validity_period {

          // group attributes:
          		:objectType = "Validity_Period" ;
          		:Validity_Start = "2007-08-13T03:33:13Z" ;
          		:Validity_Stop = "2007-08-13T05:14:37Z" ;
          } // group validity_period

        group: source {

          // group attributes:
          		:objectType = "Source" ;
          		:System = "KNMI" ;
          		:Creator = "TROPNLL2DP" ;
          		:Creator_Version = "0.9.0" ;
          		:Creation_Date = "2015-10-31T23:47:56Z" ;
          } // group source
        } // group fixed_header

      group: variable_header {

        // group attributes:
        		:objectType = "Variable_Header" ;

        group: gmd\:lineage {

          // group attributes:
          		:objectType = "gmd:LI_Lineage" ;
          		:gmd\:statement = "L2 AER_AI dataset produced by KNMI from the S5P/TROPOMI L1B product" ;

          group: gmd\:processStep {

            // group attributes:
            		:objectType = "gmi:LE_ProcessStep" ;
            		:gmd\:description = "Processing of L1b to L2 AER_AI data for orbit 4226 using the KNMI processor version 0.9.0" ;

            group: gmi\:output {

              // group attributes:
              		:objectType = "gmi:LE_Source" ;
              		:gmd\:description = "TROPOMI/S5P Aerosol Index 1-Orbit L2 Swath 7x7km" ;

              group: gmd\:sourceCitation {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;
                		:gmd\:title = "S5P_OFFL_L2__AER_AI_20070813T033313_20070813T051437_04226_01_000900_20151102T000000" ;

                group: gmd\:date {

                  // group attributes:
                  		:objectType = "gmd:CI_DateTime" ;
                  		:gmd\:date = "2015-10-31" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeListValue = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date

                group: gmd\:identifier {

                  // group attributes:
                  		:objectType = "gmd:MD_Identifier" ;
                  		:gmd\:code = "L2__AER_AI" ;
                  } // group gmd\:identifier
                } // group gmd\:sourceCitation

              group: gmi\:processedLevel {

                // group attributes:
                		:gmd\:code = "L2" ;
                		:objectType = "gmd:MD_Identifier" ;
                } // group gmi\:processedLevel
              } // group gmi\:output

            group: gmi\:processingInformation {

              // group attributes:
              		:objectType = "gmi:LE_Processing" ;

              group: gmi\:identifier {

                // group attributes:
                		:objectType = "gmd:MD_Identifier" ;
                		:gmd\:code = "KNMI L2 AER_AI processor, version 0.9.0" ;
                } // group gmi\:identifier

              group: gmi\:softwareReference {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;
                		:gmd\:title = "L2 AER_AI processor description" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "" ;
                  		:objectType = "gmd:CI_DateTime" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeListValue = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date
                } // group gmi\:softwareReference

              group: gmi\:documentation\#1 {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;
                		:gmd\:title = "TROPOMI ATBD of the UV aerosol index; S5P-KNMI-L2-0008-RP; release 1.0" ;

                group: gmd\:date {

                  // group attributes:
                  		:objectType = "gmd:CI_Date" ;
                  		:gmd\:date = "2015-11-30" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeListValue = "publication" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date
                } // group gmi\:documentation\#1

              group: gmi\:documentation\#2 {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;
                		:gmd\:title = "Sentinel-5 precursor/TROPOMI Level 2 Product User Manual UV Aerosol Index; S5P-KNMI-L2-0026-MA; release 1.0" ;

                group: gmd\:date {

                  // group attributes:
                  		:objectType = "gmd:CI_Date" ;
                  		:gmd\:date = "2015-11-30" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeListValue = "publication" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date
                } // group gmi\:documentation\#2
              } // group gmi\:processingInformation

            group: gmi\:report {

              // group attributes:
              		:gmi\:fileType = "netCDF" ;
              		:objectType = "gmi:LE_ProcessStepReport" ;
              		:gmi\:description = "Sentinel 5-precursor TROPOMI L1b processed to L2 data using the KNMI L2 AER_AI processor" ;
              		:gmi\:name = "S5P_OFFL_L2__AER_AI_20070813T033313_20070813T051437_04226_01_000900_20151102T000000.nc" ;
              } // group gmi\:report

            group: gmd\:source\#1 {

              // group attributes:
              		:objectType = "gmi:LE_Source" ;
              		:gmd\:description = "Processor CFG_AER_AI configuration file" ;

              group: gmi\:processedLevel {

                // group attributes:
                		:gmd\:code = "N/A" ;
                		:objectType = "gmd:MD_Identifier" ;
                } // group gmi\:processedLevel

              group: gmd\:sourceCitation {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2015-10-20T12:56:22Z" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeListValue = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date

                group: gmd\:title {

                  // group attributes:
                  		:gco\:characterString = "Processor CFG_AER_AI configuration file" ;
                  } // group gmd\:title

                group: gmd\:alternateTitle\#1 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_TEST_CFG_AER_AI_00000000T000000_99999999T999999_20151102T004007.cfg" ;
                  } // group gmd\:alternateTitle\#1
                } // group gmd\:sourceCitation
              } // group gmd\:source\#1

            group: gmd\:source\#2 {

              // group attributes:
              		:objectType = "gmi:LE_Source" ;
              		:gmd\:description = "TROPOMI L1B L1B_RA_BD3 radiance product" ;

              group: gmi\:processedLevel {

                // group attributes:
                		:gmd\:code = "L1B" ;
                		:objectType = "gmd:MD_Identifier" ;
                } // group gmi\:processedLevel

              group: gmd\:sourceCitation {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2015-09-30T10:22:11Z" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeListValue = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date

                group: gmd\:title {

                  // group attributes:
                  		:gco\:characterString = "TROPOMI L1B L1B_RA_BD3 radiance product" ;
                  } // group gmd\:title

                group: gmd\:alternateTitle\#1 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_TEST_L1B_RA_BD3_20070813T033313_20070813T051437_04226_02_010000_20150930T101803.nc" ;
                  } // group gmd\:alternateTitle\#1
                } // group gmd\:sourceCitation
              } // group gmd\:source\#2

            group: gmd\:source\#3 {

              // group attributes:
              		:objectType = "gmi:LE_Source" ;
              		:gmd\:description = "TROPOMI L1B L1B_IR_UVN irradiance product" ;

              group: gmi\:processedLevel {

                // group attributes:
                		:gmd\:code = "L1B" ;
                		:objectType = "gmd:MD_Identifier" ;
                } // group gmi\:processedLevel

              group: gmd\:sourceCitation {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2015-09-30T10:22:12Z" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeListValue = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date

                group: gmd\:title {

                  // group attributes:
                  		:gco\:characterString = "TROPOMI L1B L1B_IR_UVN irradiance product" ;
                  } // group gmd\:title

                group: gmd\:alternateTitle\#1 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_TEST_L1B_IR_UVN_20070813T033313_20070813T051437_04226_02_010000_20150930T101803.nc" ;
                  } // group gmd\:alternateTitle\#1
                } // group gmd\:sourceCitation
              } // group gmd\:source\#3

            group: gmd\:source\#4 {

              // group attributes:
              		:objectType = "gmi:LE_Source" ;
              		:gmd\:description = "Auxiliary ECMWF AUX_MET_2D Meteorological forecast data" ;

              group: gmi\:processedLevel {

                // group attributes:
                		:gmd\:code = "L4" ;
                		:objectType = "gmd:MD_Identifier" ;
                } // group gmi\:processedLevel

              group: gmd\:sourceCitation {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2015-05-22T08:28:55Z" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeListValue = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date

                group: gmd\:title {

                  // group attributes:
                  		:gco\:characterString = "Auxiliary ECMWF AUX_MET_2D Meteorological forecast data" ;
                  } // group gmd\:title

                group: gmd\:alternateTitle\#1 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_OFFL_AUX_MET_2D_20070812T150000_20070813T000000_20070812T120000.nc" ;
                  } // group gmd\:alternateTitle\#1

                group: gmd\:alternateTitle\#2 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_OFFL_AUX_MET_2D_20070813T030000_20070813T120000_20070813T000000.nc" ;
                  } // group gmd\:alternateTitle\#2
                } // group gmd\:sourceCitation
              } // group gmd\:source\#4

            group: gmd\:source\#5 {

              // group attributes:
              		:objectType = "gmi:LE_Source" ;
              		:gmd\:description = "Auxiliary AUX_O3___M reference data" ;

              group: gmi\:processedLevel {

                // group attributes:
                		:gmd\:code = "N/A" ;
                		:objectType = "gmd:MD_Identifier" ;
                } // group gmi\:processedLevel

              group: gmd\:sourceCitation {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2015-10-29T15:41:21Z" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeListValue = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date

                group: gmd\:title {

                  // group attributes:
                  		:gco\:characterString = "Auxiliary AUX_O3___M reference data" ;
                  } // group gmd\:title

                group: gmd\:alternateTitle\#1 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_OPER_AUX_O3___M_00000000T000000_99999999T999999_20150817T112400.nc" ;
                  } // group gmd\:alternateTitle\#1
                } // group gmd\:sourceCitation
              } // group gmd\:source\#5

            group: gmd\:source\#6 {

              // group attributes:
              		:objectType = "gmi:LE_Source" ;
              		:gmd\:description = "Auxiliary REF_DEM___ reference data" ;

              group: gmi\:processedLevel {

                // group attributes:
                		:gmd\:code = "N/A" ;
                		:objectType = "gmd:MD_Identifier" ;
                } // group gmi\:processedLevel

              group: gmd\:sourceCitation {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2015-02-06T16:58:50Z" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeListValue = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date

                group: gmd\:title {

                  // group attributes:
                  		:gco\:characterString = "Auxiliary REF_DEM___ reference data" ;
                  } // group gmd\:title

                group: gmd\:alternateTitle\#1 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_OPER_REF_DEM____00000000T000000_99999999T999999_20150206T165842.nc" ;
                  } // group gmd\:alternateTitle\#1
                } // group gmd\:sourceCitation
              } // group gmd\:source\#6

            group: gmd\:source\#7 {

              // group attributes:
              		:objectType = "gmi:LE_Source" ;
              		:gmd\:description = "Auxiliary LUT_AAI___ algorithm lookup table" ;

              group: gmi\:processedLevel {

                // group attributes:
                		:gmd\:code = "N/A" ;
                		:objectType = "gmd:MD_Identifier" ;
                } // group gmi\:processedLevel

              group: gmd\:sourceCitation {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2015-06-05T11:45:22Z" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeListValue = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date

                group: gmd\:title {

                  // group attributes:
                  		:gco\:characterString = "Auxiliary LUT_AAI___ algorithm lookup table" ;
                  } // group gmd\:title

                group: gmd\:alternateTitle\#1 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_OPER_LUT_AAI____00000000T000000_99999999T999999_20150605T114510.nc" ;
                  } // group gmd\:alternateTitle\#1
                } // group gmd\:sourceCitation
              } // group gmd\:source\#7

            group: gmd\:source\#8 {

              // group attributes:
              		:objectType = "gmi:LE_Source" ;
              		:gmd\:description = "Auxiliary REF_SOLAR_ reference data" ;

              group: gmi\:processedLevel {

                // group attributes:
                		:gmd\:code = "N/A" ;
                		:objectType = "gmd:MD_Identifier" ;
                } // group gmi\:processedLevel

              group: gmd\:sourceCitation {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2015-09-30T12:40:56Z" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeListValue = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date

                group: gmd\:title {

                  // group attributes:
                  		:gco\:characterString = "Auxiliary REF_SOLAR_ reference data" ;
                  } // group gmd\:title

                group: gmd\:alternateTitle\#1 {

                  // group attributes:
                  		:gmx\:FileName = "G2A_TEST_REF_SOLAR__00000000T000000_99999999T999999_20150930T124024.nc" ;
                  } // group gmd\:alternateTitle\#1
                } // group gmd\:sourceCitation
              } // group gmd\:source\#8

            group: gmd\:source\#9 {

              // group attributes:
              		:objectType = "gmi:LE_Source" ;
              		:gmd\:description = "Auxiliary LUT_COREG_ algorithm lookup table" ;

              group: gmi\:processedLevel {

                // group attributes:
                		:gmd\:code = "N/A" ;
                		:objectType = "gmd:MD_Identifier" ;
                } // group gmi\:processedLevel

              group: gmd\:sourceCitation {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2015-05-26T08:10:43Z" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeListValue = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date

                group: gmd\:title {

                  // group attributes:
                  		:gco\:characterString = "Auxiliary LUT_COREG_ algorithm lookup table" ;
                  } // group gmd\:title

                group: gmd\:alternateTitle\#1 {

                  // group attributes:
                  		:gmx\:FileName = "G2A_TEST_LUT_COREG__00000000T000000_99999999T999999_20150526T074640.nc" ;
                  } // group gmd\:alternateTitle\#1
                } // group gmd\:sourceCitation
              } // group gmd\:source\#9
            } // group gmd\:processStep
          } // group gmd\:lineage
        } // group variable_header
      } // group earth_explorer_header
    } // group ESA_METADATA
  } // group METADATA
}
