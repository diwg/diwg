// Contributed by Jessica Hausman <Jessica.K.Hausman AT jpl DOT nasa DOT gov>

netcdf ascat_20160616_085400_metopb_19431_eps_o_250_2401_ovw.l2 {
dimensions:
	NUMROWS = 1632 ;
	NUMCELLS = 42 ;
variables:
	int time(NUMROWS, NUMCELLS) ;
		time:_FillValue = -2147483647 ;
		time:missing_value = -2147483647 ;
		time:valid_min = 0 ;
		time:valid_max = 2147483647 ;
		time:standard_name = "time" ;
		time:long_name = "time" ;
		time:units = "seconds since 1990-01-01 00:00:00" ;
		time:coordinates = "lat lon" ;
	int lat(NUMROWS, NUMCELLS) ;
		lat:_FillValue = -2147483647 ;
		lat:missing_value = -2147483647 ;
		lat:valid_min = -9000000 ;
		lat:valid_max = 9000000 ;
		lat:standard_name = "latitude" ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:scale_factor = 1.e-05 ;
		lat:add_offset = 0. ;
	int lon(NUMROWS, NUMCELLS) ;
		lon:_FillValue = -2147483647 ;
		lon:missing_value = -2147483647 ;
		lon:valid_min = 0 ;
		lon:valid_max = 36000000 ;
		lon:standard_name = "longitude" ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:scale_factor = 1.e-05 ;
		lon:add_offset = 0. ;
	short wvc_index(NUMROWS, NUMCELLS) ;
		wvc_index:_FillValue = -32767s ;
		wvc_index:missing_value = -32767s ;
		wvc_index:valid_min = 0s ;
		wvc_index:valid_max = 999s ;
		wvc_index:standard_name = "across_swath_cell_index" ;
		wvc_index:long_name = "cross track wind vector cell number" ;
		wvc_index:units = "1" ;
		wvc_index:coordinates = "lat lon" ;
	short model_speed(NUMROWS, NUMCELLS) ;
		model_speed:_FillValue = -32767s ;
		model_speed:missing_value = -32767s ;
		model_speed:valid_min = 0s ;
		model_speed:valid_max = 5000s ;
		model_speed:standard_name = "wind_speed" ;
		model_speed:long_name = "model wind speed at 10 m" ;
		model_speed:units = "m s-1" ;
		model_speed:scale_factor = 0.01 ;
		model_speed:add_offset = 0. ;
		model_speed:coordinates = "lat lon" ;
		model_speed:background_wind_source = "ECMWF (Operational Model)" ;
	short model_dir(NUMROWS, NUMCELLS) ;
		model_dir:_FillValue = -32767s ;
		model_dir:missing_value = -32767s ;
		model_dir:valid_min = 0s ;
		model_dir:valid_max = 3600s ;
		model_dir:standard_name = "wind_to_direction" ;
		model_dir:long_name = "model wind direction at 10 m" ;
		model_dir:units = "degree" ;
		model_dir:scale_factor = 0.1 ;
		model_dir:add_offset = 0. ;
		model_dir:coordinates = "lat lon" ;
		model_dir:background_wind_source = "ECMWF (Operational Model)" ;
	short ice_prob(NUMROWS, NUMCELLS) ;
		ice_prob:_FillValue = -32767s ;
		ice_prob:missing_value = -32767s ;
		ice_prob:valid_min = 0s ;
		ice_prob:valid_max = 1000s ;
		ice_prob:long_name = "ice probability" ;
		ice_prob:units = "1" ;
		ice_prob:scale_factor = 0.001 ;
		ice_prob:add_offset = 0. ;
		ice_prob:coordinates = "lat lon" ;
	short ice_age(NUMROWS, NUMCELLS) ;
		ice_age:_FillValue = -32767s ;
		ice_age:missing_value = -32767s ;
		ice_age:valid_min = -5000s ;
		ice_age:valid_max = 5000s ;
		ice_age:long_name = "ice age (a-parameter)" ;
		ice_age:units = "dB" ;
		ice_age:scale_factor = 0.01 ;
		ice_age:add_offset = 0. ;
		ice_age:coordinates = "lat lon" ;
	int wvc_quality_flag(NUMROWS, NUMCELLS) ;
		wvc_quality_flag:_FillValue = -2147483647 ;
		wvc_quality_flag:missing_value = -2147483647 ;
		wvc_quality_flag:valid_min = 0 ;
		wvc_quality_flag:valid_max = 8388607 ;
		wvc_quality_flag:standard_name = "status_flag" ;
		wvc_quality_flag:long_name = "wind vector cell quality" ;
		wvc_quality_flag:coordinates = "lat lon" ;
		wvc_quality_flag:flag_masks = 64, 128, 256, 512, 1024, 2048, 4096, 8192, 16384, 32768, 65536, 131072, 262144, 524288, 1048576, 2097152, 4194304 ;
		wvc_quality_flag:flag_meanings = "distance_to_gmf_too_large data_are_redundant no_meteorological_background_used rain_detected rain_flag_not_usable small_wind_less_than_or_equal_to_3_m_s large_wind_greater_than_30_m_s wind_inversion_not_successful some_portion_of_wvc_is_over_ice some_portion_of_wvc_is_over_land variational_quality_control_fails knmi_quality_control_fails product_monitoring_event_flag product_monitoring_not_used any_beam_noise_content_above_threshold poor_azimuth_diversity not_enough_good_sigma0_for_wind_retrieval" ;
	short wind_speed(NUMROWS, NUMCELLS) ;
		wind_speed:_FillValue = -32767s ;
		wind_speed:missing_value = -32767s ;
		wind_speed:valid_min = 0s ;
		wind_speed:valid_max = 5000s ;
		wind_speed:standard_name = "wind_speed" ;
		wind_speed:long_name = "wind speed at 10 m" ;
		wind_speed:units = "m s-1" ;
		wind_speed:scale_factor = 0.01 ;
		wind_speed:add_offset = 0. ;
		wind_speed:coordinates = "lat lon" ;
	short wind_dir(NUMROWS, NUMCELLS) ;
		wind_dir:_FillValue = -32767s ;
		wind_dir:missing_value = -32767s ;
		wind_dir:valid_min = 0s ;
		wind_dir:valid_max = 3600s ;
		wind_dir:standard_name = "wind_to_direction" ;
		wind_dir:long_name = "wind direction at 10 m" ;
		wind_dir:units = "degree" ;
		wind_dir:scale_factor = 0.1 ;
		wind_dir:add_offset = 0. ;
		wind_dir:coordinates = "lat lon" ;
	short bs_distance(NUMROWS, NUMCELLS) ;
		bs_distance:_FillValue = -32767s ;
		bs_distance:missing_value = -32767s ;
		bs_distance:valid_min = -500s ;
		bs_distance:valid_max = 500s ;
		bs_distance:standard_name = "backscatter_distance_to_modelfunction" ;
		bs_distance:long_name = "backscatter distance" ;
		bs_distance:units = "1" ;
		bs_distance:scale_factor = 0.1 ;
		bs_distance:add_offset = 0. ;
		bs_distance:coordinates = "lat lon" ;

// global attributes:
		:title = "MetOp-B ASCAT Level 2 25.0 km Ocean Surface Wind Vector Product" ;
		:title_short_name = "ASCATB-L2-25km" ;
		:Conventions = "CF-1.4" ;
		:institution = "EUMETSAT/OSI SAF/KNMI" ;
		:source = "MetOp-B ASCAT" ;
		:software_identification_level_1 = 1000 ;
		:instrument_calibration_version = 0 ;
		:software_identification_wind = 2401 ;
		:pixel_size_on_horizontal = "25.0 km" ;
		:service_type = "eps" ;
		:processing_type = "O" ;
		:contents = "ovw" ;
		:granule_name = "ascat_20160616_085400_metopb_19431_eps_o_250_2401_ovw.l2.nc" ;
		:processing_level = "L2" ;
		:orbit_number = 19431 ;
		:start_date = "2016-06-16" ;
		:start_time = "08:54:00" ;
		:stop_date = "2016-06-16" ;
		:stop_time = "10:35:56" ;
		:equator_crossing_longitude = " 189.571" ;
		:equator_crossing_date = "2016-06-16" ;
		:equator_crossing_time = "08:51:59" ;
		:rev_orbit_period = "6081.7" ;
		:orbit_inclination = "98.7" ;
		:history = "N/A" ;
		:references = "ASCAT Wind Product User Manual, http://www.osi-saf.org/, http://www.knmi.nl/scatterometer/" ;
		:comment = "Orbit period and inclination are constant values. All wind directions in oceanographic convention (0 deg. flowing North)" ;
		:creation_date = "2016-06-16" ;
		:creation_time = "11:26:13" ;
}
