// -*-C++-*-

// Purpose: CDL file to demonstrate best practices for curvilinear datasets, aka, Swaths
// Part of an ongoing project by NASA's Dataset Interoperability Working Group (DIWG)
// Comments, questions, suggestions to fxm

// Usage:
// ncgen             -b -o swath_modis_l2.nc swath_modis_l2.cdl # netCDF3
// ncgen -k netCDF-4 -b -o swath_modis_l2.nc swath_modis_l2.cdl # netCDF4

// URL: 
// git clone http://github.com/diwg/diwg.git
// http://github.com/diwg/diwg/swath_modis_l2.cdl

netcdf swath_modis_l2 {

// Template source: MOD04_L2.A2010091.0950.051.2010104212718.hdf
  dimensions:
    Xtrack = 3 ;
    Track = 2 ;
    Band = 2 ;

  variables:
    double Band(Band) ;
      Band:long_name = "Wavelength" ;
      Band:units = "micron" ;

    double Latitude(Track,Xtrack) ;
      Latitude:long_name = "Geodetic Latitude" ;
      Latitude:units = "Degrees_north" ;
      Latitude:Track_Sampling = 5, 2025, 10 ;
      Latitude:Xtrack_Sampling = 5, 1345, 10 ;
      Latitude:Geolocation_Pointer = "Geolocation data not applicable" ;

    double Longitude(Track,Xtrack) ;
      Longitude:long_name = "Geodetic Longitude" ;
      Longitude:units = "Degrees_east" ;
      Longitude:Track_Sampling = 5, 2025, 10 ;
      Longitude:Xtrack_Sampling = 5, 1345, 10 ;
      Longitude:Geolocation_Pointer = "Geolocation data not applicable" ;

    short AOD550(Track,Xtrack) ;
      AOD550:valid_range = 0s, 5000s ;
      AOD550:_FillValue = -9999s ;
      AOD550:long_name = "AOT at 0.55 micron" ;
      AOD550:units = "None" ;
      AOD550:scale_factor = 0.001f ;
      AOD550:add_offset = 0.0f ;
      AOD550:Track_Sampling = 5, 2025, 10 ;
      AOD550:Xtrack_Sampling = 5, 1345, 10 ;
      AOD550:Geolocation_Pointer = "Internal geolocation arrays" ;

    short AOD_spectral(Band,Track,Xtrack) ;
      AOD_spectral:valid_range = -100s, 5000s ;
      AOD_spectral:_FillValue = -9999s ;
      AOD_spectral:long_name = "AOT every band" ;
      AOD_spectral:units = "None" ;
      AOD_spectral:scale_factor = 0.001f ;
      AOD_spectral:add_offset = 0.0f ;

      data:
	Band=500,550;
	Latitude=-45,-44,-43,45,46,47;
	Longitude=-120,-119,0,1,120,121;
	AOD550=1,2,3,4,5,6;
	AOD_spectral=1,2,3,4,5,6,7,8,9,10,11,12;
} // group /
