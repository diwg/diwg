netcdf S5P_TEST_L1B_IR_UVN_20140827T114200_20140827T115800_53811_01_000901_20141209T120000 {

// global attributes:
		:time_coverage_end = "2014-08-27T11:52:00Z" ;
		:time_coverage_start = "2014-08-27T11:51:48Z" ;
		:time_reference = "2014-08-27T00:00:00Z" ;

group: BAND1_IRRADIANCE {

  group: STANDARD_MODE {
    dimensions:
    	time = 1 ;
    	pixel = 76 ;
    	spectral_channel = 497 ;
    	scanline = 1 ;
    	nsettings = 1 ;
    	nbinningregions = 18 ;

    group: OBSERVATIONS {
      variables:
      	int pixel(pixel) ;
      		pixel:comment = "This dimension variable defines the indices across track; index starts at 0" ;
      		pixel:long_name = "across track dimension index" ;
      		pixel:units = "1" ;
      	int spectral_channel(spectral_channel) ;
      		spectral_channel:comment = "This dimension variable defines the indices spectral dimension; index starts at 0" ;
      		spectral_channel:long_name = "wavelength dimension index" ;
      		spectral_channel:units = "1" ;
      	int scanline(scanline) ;
      		scanline:comment = "This dimension variable defines the indices along track; index starts at 0" ;
      		scanline:long_name = "along track dimension index" ;
      		scanline:units = "1" ;
      	int delta_time(time, scanline) ;
      		delta_time:comment = "Time difference with time for each measurement" ;
      		delta_time:_FillValue = -2147483647 ;
      		delta_time:long_name = "offset from the reference start time of measurement" ;
      		delta_time:units = "milliseconds since 2014-08-27 00:00:00" ;
      	ushort detector_column_qualification(time, scanline, spectral_channel) ;
      		detector_column_qualification:comment = "Qualification flag indicating column indicating column type or state" ;
      		detector_column_qualification:_FillValue = 65535US ;
      		detector_column_qualification:flag_values = 0US, 1US, 16US, 32US, 64US, 256US, 512US, 1024US, 2048US ;
      		detector_column_qualification:flag_masks = 0US, 1US, 16US, 98US, 98US, 3840US, 3840US, 3840US, 3840US ;
      		detector_column_qualification:flag_meanings = "no_qualification skipped uvn_odd uvn_prepost uvn_overscan swir_adc0 swir_adc1 swir_adc2 swir_adc3" ;
      		detector_column_qualification:long_name = "Detector column qualification flags" ;
      		detector_column_qualification:max_val = 65534US ;
      		detector_column_qualification:min_val = 0US ;
      		detector_column_qualification:units = "1" ;
      	ushort detector_row_qualification(time, scanline, pixel) ;
      		detector_row_qualification:comment = "Qualification flag indicating row type or state" ;
      		detector_row_qualification:_FillValue = 65535US ;
      		detector_row_qualification:flag_values = 0US, 1US, 2US, 4US, 8US, 16US, 256US, 4096US, 8192US ;
      		detector_row_qualification:flag_masks = 0US, 9US, 2US, 4US, 9US, 16US, 256US, 4096US, 8192US ;
      		detector_row_qualification:flag_meanings = "no_qualification uvn_ror uvn_dump uvn_covered uvn_overscan uvn_higain swir_reference gen_transistion gen_non_illuminated" ;
      		detector_row_qualification:long_name = "Detector row qualification flags" ;
      		detector_row_qualification:max_val = 65534US ;
      		detector_row_qualification:min_val = 0US ;
      		detector_row_qualification:units = "1" ;
      	ushort measurement_quality(time, scanline) ;
      		measurement_quality:flag_values = 0US, 1US, 2US, 16US, 32US, 128US, 256US, 4096US ;
      		measurement_quality:flag_masks = 0US, 1US, 2US, 16US, 32US, 128US, 256US, 4096US ;
      		measurement_quality:flag_meanings = "no_error proc_skipped no_residual saa spacecraft_manoeuvre sub_grp irr_out_of_range sub_group" ;
      		measurement_quality:long_name = "measurement quality flag" ;
      		measurement_quality:max_val = 65534US ;
      		measurement_quality:min_val = 0US ;
      		measurement_quality:units = "1" ;
      		measurement_quality:comment = "Overall quality information for a measurement" ;
      		measurement_quality:coordinates = "longitude latitude" ;
      		measurement_quality:_FillValue = 65535US ;
      	float irradiance(time, scanline, pixel, spectral_channel) ;
      		irradiance:ancilary_vars = "irradiance_noise irradiance_error quality_level spectral_channel_quality" ;
      		irradiance:comment = "Measured spectral irradiance for each spectral pixel" ;
      		irradiance:_FillValue = 9.96921e+36f ;
      		irradiance:long_name = "spectral photon irradiance" ;
      		irradiance:units = "mol.m-2.nm-1.s-1" ;
      	byte irradiance_error(time, scanline, pixel, spectral_channel) ;
      		irradiance_error:comment = "The irradiance_error is a measure for the one standard deviation error of the bias of the irradiance measurement; it is expressed in decibel (dB), i.e. 10 times the base-10 logarithmic value of the ratio between the irradiance and the estimation error." ;
      		irradiance_error:coordinates = "longitude latitude" ;
      		irradiance_error:_FillValue = -127b ;
      		irradiance_error:long_name = "spectral irradiance noise" ;
      		irradiance_error:units = "1" ;
      	byte irradiance_noise(time, scanline, pixel, spectral_channel) ;
      		irradiance_noise:comment = "The irradiance_noise is a measure for the one standard deviation random error of the irradiance measurement; it is expressed in decibel (dB), i.e. 10 times the base-10 logarithmic value of the ratio between the irradiance and the random error." ;
      		irradiance_noise:coordinates = "longitude latitude" ;
      		irradiance_noise:_FillValue = -127b ;
      		irradiance_noise:long_name = "spectral photon irradiance noise, one standard deviation" ;
      		irradiance_noise:units = "1" ;
      	ubyte quality_level(time, scanline, pixel, spectral_channel) ;
      		quality_level:comment = "Overall quality assessment information for each (spectral) pixel" ;
      		quality_level:coordinates = "longitude latitude" ;
      		quality_level:_FillValue = 255UB ;
      		quality_level:long_name = "qualiy level of spectral channel" ;
      		quality_level:max_val = 100UB ;
      		quality_level:min_val = 0UB ;
      		quality_level:units = "mol.m-2.nm-1.s-1" ;
      	ubyte spectral_channel_quality(time, scanline, pixel, spectral_channel) ;
      		spectral_channel_quality:comment = "Quality assessment information for each (spectral) pixel" ;
      		spectral_channel_quality:coordinates = "longitude latitude" ;
      		spectral_channel_quality:_FillValue = 255UB ;
      		spectral_channel_quality:flag_values = 0UB, 1UB, 2UB, 8UB, 16UB, 32UB, 64UB, 128UB ;
      		spectral_channel_quality:flag_masks = 0UB, 1UB, 2UB, 8UB, 16UB, 32UB, 64UB, 128UB ;
      		spectral_channel_quality:flag_meanings = "no_error missing bad_pixel processing_error saturated transient rts underflow" ;
      		spectral_channel_quality:long_name = "spectral channel quality flag" ;
      		spectral_channel_quality:max_val = 254UB ;
      		spectral_channel_quality:min_val = 0UB ;
      		spectral_channel_quality:units = "mol.m-2.nm-1.s-1" ;
      	int time(time) ;
      		time:comment = "Reference time of the measurements. The reference time is set to yyyy-mm-ddT00:00:00 UTC, where yyyy-mm-dd is the day on which the measurements of a particular data granule start." ;
      		time:long_name = "reference start time of measurement" ;
      		time:standard_name = "time" ;
      		time:units = "seconds since 2010-01-01 00:00:00" ;
      } // group OBSERVATIONS

    group: GEODATA {
      variables:
      	float earth_sun_distance(time) ;
      		earth_sun_distance:comment = "1 ua equals 149,597,870,700 meters" ;
      		earth_sun_distance:_FillValue = 9.96921e+36f ;
      		earth_sun_distance:long_name = "distance between the earth and the sun" ;
      		earth_sun_distance:max_val = 1.02f ;
      		earth_sun_distance:min_val = 0.98f ;
      		earth_sun_distance:units = "ua" ;
      } // group GEODATA
    } // group STANDARD_MODE
  } // group BAND1_IRRADIANCE

group: BAND2_IRRADIANCE {

  group: STANDARD_MODE {
    dimensions:
    	time = 1 ;
    	pixel = 308 ;
    	spectral_channel = 497 ;
    	scanline = 1 ;
    	nsettings = 1 ;
    	nbinningregions = 18 ;

    group: OBSERVATIONS {
      variables:
      	int pixel(pixel) ;
      		pixel:comment = "This dimension variable defines the indices across track; index starts at 0" ;
      		pixel:long_name = "across track dimension index" ;
      		pixel:units = "1" ;
      	int spectral_channel(spectral_channel) ;
      		spectral_channel:comment = "This dimension variable defines the indices spectral dimension; index starts at 0" ;
      		spectral_channel:long_name = "wavelength dimension index" ;
      		spectral_channel:units = "1" ;
      	int scanline(scanline) ;
      		scanline:comment = "This dimension variable defines the indices along track; index starts at 0" ;
      		scanline:long_name = "along track dimension index" ;
      		scanline:units = "1" ;
      	int delta_time(time, scanline) ;
      		delta_time:comment = "Time difference with time for each measurement" ;
      		delta_time:_FillValue = -2147483647 ;
      		delta_time:long_name = "offset from the reference start time of measurement" ;
      		delta_time:units = "milliseconds since 2014-08-27 00:00:00" ;
      	ushort detector_column_qualification(time, scanline, spectral_channel) ;
      		detector_column_qualification:comment = "Qualification flag indicating column indicating column type or state" ;
      		detector_column_qualification:_FillValue = 65535US ;
      		detector_column_qualification:flag_values = 0US, 1US, 16US, 32US, 64US, 256US, 512US, 1024US, 2048US ;
      		detector_column_qualification:flag_masks = 0US, 1US, 16US, 98US, 98US, 3840US, 3840US, 3840US, 3840US ;
      		detector_column_qualification:flag_meanings = "no_qualification skipped uvn_odd uvn_prepost uvn_overscan swir_adc0 swir_adc1 swir_adc2 swir_adc3" ;
      		detector_column_qualification:long_name = "Detector column qualification flags" ;
      		detector_column_qualification:max_val = 65534US ;
      		detector_column_qualification:min_val = 0US ;
      		detector_column_qualification:units = "1" ;
      	ushort detector_row_qualification(time, scanline, pixel) ;
      		detector_row_qualification:comment = "Qualification flag indicating row type or state" ;
      		detector_row_qualification:_FillValue = 65535US ;
      		detector_row_qualification:flag_values = 0US, 1US, 2US, 4US, 8US, 16US, 256US, 4096US, 8192US ;
      		detector_row_qualification:flag_masks = 0US, 9US, 2US, 4US, 9US, 16US, 256US, 4096US, 8192US ;
      		detector_row_qualification:flag_meanings = "no_qualification uvn_ror uvn_dump uvn_covered uvn_overscan uvn_higain swir_reference gen_transistion gen_non_illuminated" ;
      		detector_row_qualification:long_name = "Detector row qualification flags" ;
      		detector_row_qualification:max_val = 65534US ;
      		detector_row_qualification:min_val = 0US ;
      		detector_row_qualification:units = "1" ;
      	ushort measurement_quality(time, scanline) ;
      		measurement_quality:flag_values = 0US, 1US, 2US, 16US, 32US, 128US, 256US, 4096US ;
      		measurement_quality:flag_masks = 0US, 1US, 2US, 16US, 32US, 128US, 256US, 4096US ;
      		measurement_quality:flag_meanings = "no_error proc_skipped no_residual saa spacecraft_manoeuvre sub_grp irr_out_of_range sub_group" ;
      		measurement_quality:long_name = "measurement quality flag" ;
      		measurement_quality:max_val = 65534US ;
      		measurement_quality:min_val = 0US ;
      		measurement_quality:units = "1" ;
      		measurement_quality:comment = "Overall quality information for a measurement" ;
      		measurement_quality:coordinates = "longitude latitude" ;
      		measurement_quality:_FillValue = 65535US ;
      	float irradiance(time, scanline, pixel, spectral_channel) ;
      		irradiance:ancilary_vars = "irradiance_noise irradiance_error quality_level spectral_channel_quality" ;
      		irradiance:comment = "Measured spectral irradiance for each spectral pixel" ;
      		irradiance:_FillValue = 9.96921e+36f ;
      		irradiance:long_name = "spectral photon irradiance" ;
      		irradiance:units = "mol.m-2.nm-1.s-1" ;
      	byte irradiance_error(time, scanline, pixel, spectral_channel) ;
      		irradiance_error:comment = "The irradiance_error is a measure for the one standard deviation error of the bias of the irradiance measurement; it is expressed in decibel (dB), i.e. 10 times the base-10 logarithmic value of the ratio between the irradiance and the estimation error." ;
      		irradiance_error:units = "1" ;
      		irradiance_error:coordinates = "longitude latitude" ;
      		irradiance_error:_FillValue = -127b ;
      		irradiance_error:long_name = "spectral irradiance noise" ;
      	byte irradiance_noise(time, scanline, pixel, spectral_channel) ;
      		irradiance_noise:comment = "The irradiance_noise is a measure for the one standard deviation random error of the irradiance measurement; it is expressed in decibel (dB), i.e. 10 times the base-10 logarithmic value of the ratio between the irradiance and the random error." ;
      		irradiance_noise:coordinates = "longitude latitude" ;
      		irradiance_noise:_FillValue = -127b ;
      		irradiance_noise:long_name = "spectral photon irradiance noise, one standard deviation" ;
      		irradiance_noise:units = "1" ;
      	ubyte quality_level(time, scanline, pixel, spectral_channel) ;
      		quality_level:comment = "Overall quality assessment information for each (spectral) pixel" ;
      		quality_level:coordinates = "longitude latitude" ;
      		quality_level:_FillValue = 255UB ;
      		quality_level:long_name = "qualiy level of spectral channel" ;
      		quality_level:max_val = 100UB ;
      		quality_level:min_val = 0UB ;
      		quality_level:units = "mol.m-2.nm-1.s-1" ;
      	ubyte spectral_channel_quality(time, scanline, pixel, spectral_channel) ;
      		spectral_channel_quality:comment = "Quality assessment information for each (spectral) pixel" ;
      		spectral_channel_quality:coordinates = "longitude latitude" ;
      		spectral_channel_quality:_FillValue = 255UB ;
      		spectral_channel_quality:max_val = 254UB ;
      		spectral_channel_quality:flag_values = 0UB, 1UB, 2UB, 8UB, 16UB, 32UB, 64UB, 128UB ;
      		spectral_channel_quality:flag_masks = 0UB, 1UB, 2UB, 8UB, 16UB, 32UB, 64UB, 128UB ;
      		spectral_channel_quality:flag_meanings = "no_error missing bad_pixel processing_error saturated transient rts underflow" ;
      		spectral_channel_quality:long_name = "spectral channel quality flag" ;
      		spectral_channel_quality:min_val = 0UB ;
      		spectral_channel_quality:units = "mol.m-2.nm-1.s-1" ;
      	int time(time) ;
      		time:comment = "Reference time of the measurements. The reference time is set to yyyy-mm-ddT00:00:00 UTC, where yyyy-mm-dd is the day on which the measurements of a particular data granule start." ;
      		time:long_name = "reference start time of measurement" ;
      		time:standard_name = "time" ;
      		time:units = "seconds since 2010-01-01 00:00:00" ;
      } // group OBSERVATIONS

    group: GEODATA {
      variables:
      	float earth_sun_distance(time) ;
      		earth_sun_distance:comment = "1 ua equals 149,597,870,700 meters" ;
      		earth_sun_distance:_FillValue = 9.96921e+36f ;
      		earth_sun_distance:long_name = "distance between the earth and the sun" ;
      		earth_sun_distance:max_val = 1.02f ;
      		earth_sun_distance:min_val = 0.98f ;
      		earth_sun_distance:units = "ua" ;
      } // group GEODATA
    } // group STANDARD_MODE
  } // group BAND2_IRRADIANCE

group: BAND3_IRRADIANCE {

  group: STANDARD_MODE {
    dimensions:
    	time = 1 ;
    	pixel = 309 ;
    	spectral_channel = 497 ;
    	scanline = 1 ;
    	nsettings = 1 ;
    	nbinningregions = 18 ;

    group: OBSERVATIONS {
      variables:
      	int pixel(pixel) ;
      		pixel:comment = "This dimension variable defines the indices across track; index starts at 0" ;
      		pixel:long_name = "across track dimension index" ;
      		pixel:units = "1" ;
      	int spectral_channel(spectral_channel) ;
      		spectral_channel:comment = "This dimension variable defines the indices spectral dimension; index starts at 0" ;
      		spectral_channel:long_name = "wavelength dimension index" ;
      		spectral_channel:units = "1" ;
      	int scanline(scanline) ;
      		scanline:comment = "This dimension variable defines the indices along track; index starts at 0" ;
      		scanline:long_name = "along track dimension index" ;
      		scanline:units = "1" ;
      	int delta_time(time, scanline) ;
      		delta_time:comment = "Time difference with time for each measurement" ;
      		delta_time:_FillValue = -2147483647 ;
      		delta_time:long_name = "offset from the reference start time of measurement" ;
      		delta_time:units = "milliseconds since 2014-08-27 00:00:00" ;
      	ushort detector_column_qualification(time, scanline, spectral_channel) ;
      		detector_column_qualification:comment = "Qualification flag indicating column indicating column type or state" ;
      		detector_column_qualification:_FillValue = 65535US ;
      		detector_column_qualification:flag_values = 0US, 1US, 16US, 32US, 64US, 256US, 512US, 1024US, 2048US ;
      		detector_column_qualification:flag_masks = 0US, 1US, 16US, 98US, 98US, 3840US, 3840US, 3840US, 3840US ;
      		detector_column_qualification:flag_meanings = "no_qualification skipped uvn_odd uvn_prepost uvn_overscan swir_adc0 swir_adc1 swir_adc2 swir_adc3" ;
      		detector_column_qualification:long_name = "Detector column qualification flags" ;
      		detector_column_qualification:max_val = 65534US ;
      		detector_column_qualification:min_val = 0US ;
      		detector_column_qualification:units = "1" ;
      	ushort detector_row_qualification(time, scanline, pixel) ;
      		detector_row_qualification:comment = "Qualification flag indicating row type or state" ;
      		detector_row_qualification:_FillValue = 65535US ;
      		detector_row_qualification:flag_values = 0US, 1US, 2US, 4US, 8US, 16US, 256US, 4096US, 8192US ;
      		detector_row_qualification:flag_masks = 0US, 9US, 2US, 4US, 9US, 16US, 256US, 4096US, 8192US ;
      		detector_row_qualification:flag_meanings = "no_qualification uvn_ror uvn_dump uvn_covered uvn_overscan uvn_higain swir_reference gen_transistion gen_non_illuminated" ;
      		detector_row_qualification:long_name = "Detector row qualification flags" ;
      		detector_row_qualification:max_val = 65534US ;
      		detector_row_qualification:min_val = 0US ;
      		detector_row_qualification:units = "1" ;
      	ushort measurement_quality(time, scanline) ;
      		measurement_quality:flag_values = 0US, 1US, 2US, 16US, 32US, 128US, 256US, 4096US ;
      		measurement_quality:flag_masks = 0US, 1US, 2US, 16US, 32US, 128US, 256US, 4096US ;
      		measurement_quality:flag_meanings = "no_error proc_skipped no_residual saa spacecraft_manoeuvre sub_grp irr_out_of_range sub_group" ;
      		measurement_quality:long_name = "measurement quality flag" ;
      		measurement_quality:max_val = 65534US ;
      		measurement_quality:min_val = 0US ;
      		measurement_quality:units = "1" ;
      		measurement_quality:comment = "Overall quality information for a measurement" ;
      		measurement_quality:coordinates = "longitude latitude" ;
      		measurement_quality:_FillValue = 65535US ;
      	float irradiance(time, scanline, pixel, spectral_channel) ;
      		irradiance:ancilary_vars = "irradiance_noise irradiance_error quality_level spectral_channel_quality" ;
      		irradiance:comment = "Measured spectral irradiance for each spectral pixel" ;
      		irradiance:long_name = "spectral photon irradiance" ;
      		irradiance:_FillValue = 9.96921e+36f ;
      		irradiance:units = "mol.m-2.nm-1.s-1" ;
      	byte irradiance_error(time, scanline, pixel, spectral_channel) ;
      		irradiance_error:comment = "The irradiance_error is a measure for the one standard deviation error of the bias of the irradiance measurement; it is expressed in decibel (dB), i.e. 10 times the base-10 logarithmic value of the ratio between the irradiance and the estimation error." ;
      		irradiance_error:coordinates = "longitude latitude" ;
      		irradiance_error:_FillValue = -127b ;
      		irradiance_error:long_name = "spectral irradiance noise" ;
      		irradiance_error:units = "1" ;
      	byte irradiance_noise(time, scanline, pixel, spectral_channel) ;
      		irradiance_noise:comment = "The irradiance_noise is a measure for the one standard deviation random error of the irradiance measurement; it is expressed in decibel (dB), i.e. 10 times the base-10 logarithmic value of the ratio between the irradiance and the random error." ;
      		irradiance_noise:coordinates = "longitude latitude" ;
      		irradiance_noise:_FillValue = -127b ;
      		irradiance_noise:long_name = "spectral photon irradiance noise, one standard deviation" ;
      		irradiance_noise:units = "1" ;
      	ubyte quality_level(time, scanline, pixel, spectral_channel) ;
      		quality_level:comment = "Overall quality assessment information for each (spectral) pixel" ;
      		quality_level:coordinates = "longitude latitude" ;
      		quality_level:_FillValue = 255UB ;
      		quality_level:long_name = "qualiy level of spectral channel" ;
      		quality_level:max_val = 100UB ;
      		quality_level:min_val = 0UB ;
      		quality_level:units = "mol.m-2.nm-1.s-1" ;
      	ubyte spectral_channel_quality(time, scanline, pixel, spectral_channel) ;
      		spectral_channel_quality:comment = "Quality assessment information for each (spectral) pixel" ;
      		spectral_channel_quality:coordinates = "longitude latitude" ;
      		spectral_channel_quality:_FillValue = 255UB ;
      		spectral_channel_quality:flag_values = 0UB, 1UB, 2UB, 8UB, 16UB, 32UB, 64UB, 128UB ;
      		spectral_channel_quality:flag_masks = 0UB, 1UB, 2UB, 8UB, 16UB, 32UB, 64UB, 128UB ;
      		spectral_channel_quality:flag_meanings = "no_error missing bad_pixel processing_error saturated transient rts underflow" ;
      		spectral_channel_quality:long_name = "spectral channel quality flag" ;
      		spectral_channel_quality:max_val = 254UB ;
      		spectral_channel_quality:min_val = 0UB ;
      		spectral_channel_quality:units = "mol.m-2.nm-1.s-1" ;
      	int time(time) ;
      		time:comment = "Reference time of the measurements. The reference time is set to yyyy-mm-ddT00:00:00 UTC, where yyyy-mm-dd is the day on which the measurements of a particular data granule start." ;
      		time:long_name = "reference start time of measurement" ;
      		time:standard_name = "time" ;
      		time:units = "seconds since 2010-01-01 00:00:00" ;
      } // group OBSERVATIONS

    group: GEODATA {
      variables:
      	float earth_sun_distance(time) ;
      		earth_sun_distance:comment = "1 ua equals 149,597,870,700 meters" ;
      		earth_sun_distance:_FillValue = 9.96921e+36f ;
      		earth_sun_distance:long_name = "distance between the earth and the sun" ;
      		earth_sun_distance:max_val = 1.02f ;
      		earth_sun_distance:min_val = 0.98f ;
      		earth_sun_distance:units = "ua" ;
      } // group GEODATA
    } // group STANDARD_MODE
  } // group BAND3_IRRADIANCE

group: BAND4_IRRADIANCE {

  group: STANDARD_MODE {
    dimensions:
    	time = 1 ;
    	pixel = 309 ;
    	spectral_channel = 497 ;
    	scanline = 1 ;
    	nsettings = 1 ;
    	nbinningregions = 18 ;

    group: OBSERVATIONS {
      variables:
      	int pixel(pixel) ;
      		pixel:comment = "This dimension variable defines the indices across track; index starts at 0" ;
      		pixel:long_name = "across track dimension index" ;
      		pixel:units = "1" ;
      	int spectral_channel(spectral_channel) ;
      		spectral_channel:comment = "This dimension variable defines the indices spectral dimension; index starts at 0" ;
      		spectral_channel:long_name = "wavelength dimension index" ;
      		spectral_channel:units = "1" ;
      	int scanline(scanline) ;
      		scanline:comment = "This dimension variable defines the indices along track; index starts at 0" ;
      		scanline:long_name = "along track dimension index" ;
      		scanline:units = "1" ;
      	int delta_time(time, scanline) ;
      		delta_time:comment = "Time difference with time for each measurement" ;
      		delta_time:_FillValue = -2147483647 ;
      		delta_time:long_name = "offset from the reference start time of measurement" ;
      		delta_time:units = "milliseconds since 2014-08-27 00:00:00" ;
      	ushort detector_column_qualification(time, scanline, spectral_channel) ;
      		detector_column_qualification:comment = "Qualification flag indicating column indicating column type or state" ;
      		detector_column_qualification:_FillValue = 65535US ;
      		detector_column_qualification:flag_values = 0US, 1US, 16US, 32US, 64US, 256US, 512US, 1024US, 2048US ;
      		detector_column_qualification:flag_masks = 0US, 1US, 16US, 98US, 98US, 3840US, 3840US, 3840US, 3840US ;
      		detector_column_qualification:flag_meanings = "no_qualification skipped uvn_odd uvn_prepost uvn_overscan swir_adc0 swir_adc1 swir_adc2 swir_adc3" ;
      		detector_column_qualification:long_name = "Detector column qualification flags" ;
      		detector_column_qualification:max_val = 65534US ;
      		detector_column_qualification:min_val = 0US ;
      		detector_column_qualification:units = "1" ;
      	ushort detector_row_qualification(time, scanline, pixel) ;
      		detector_row_qualification:comment = "Qualification flag indicating row type or state" ;
      		detector_row_qualification:_FillValue = 65535US ;
      		detector_row_qualification:flag_values = 0US, 1US, 2US, 4US, 8US, 16US, 256US, 4096US, 8192US ;
      		detector_row_qualification:flag_masks = 0US, 9US, 2US, 4US, 9US, 16US, 256US, 4096US, 8192US ;
      		detector_row_qualification:flag_meanings = "no_qualification uvn_ror uvn_dump uvn_covered uvn_overscan uvn_higain swir_reference gen_transistion gen_non_illuminated" ;
      		detector_row_qualification:long_name = "Detector row qualification flags" ;
      		detector_row_qualification:max_val = 65534US ;
      		detector_row_qualification:min_val = 0US ;
      		detector_row_qualification:units = "1" ;
      	ushort measurement_quality(time, scanline) ;
      		measurement_quality:flag_values = 0US, 1US, 2US, 16US, 32US, 128US, 256US, 4096US ;
      		measurement_quality:flag_masks = 0US, 1US, 2US, 16US, 32US, 128US, 256US, 4096US ;
      		measurement_quality:flag_meanings = "no_error proc_skipped no_residual saa spacecraft_manoeuvre sub_grp irr_out_of_range sub_group" ;
      		measurement_quality:long_name = "measurement quality flag" ;
      		measurement_quality:max_val = 65534US ;
      		measurement_quality:min_val = 0US ;
      		measurement_quality:units = "1" ;
      		measurement_quality:comment = "Overall quality information for a measurement" ;
      		measurement_quality:coordinates = "longitude latitude" ;
      		measurement_quality:_FillValue = 65535US ;
      	float irradiance(time, scanline, pixel, spectral_channel) ;
      		irradiance:ancilary_vars = "irradiance_noise irradiance_error quality_level spectral_channel_quality" ;
      		irradiance:comment = "Measured spectral irradiance for each spectral pixel" ;
      		irradiance:units = "mol.m-2.nm-1.s-1" ;
      		irradiance:_FillValue = 9.96921e+36f ;
      		irradiance:long_name = "spectral photon irradiance" ;
      	byte irradiance_error(time, scanline, pixel, spectral_channel) ;
      		irradiance_error:comment = "The irradiance_error is a measure for the one standard deviation error of the bias of the irradiance measurement; it is expressed in decibel (dB), i.e. 10 times the base-10 logarithmic value of the ratio between the irradiance and the estimation error." ;
      		irradiance_error:coordinates = "longitude latitude" ;
      		irradiance_error:_FillValue = -127b ;
      		irradiance_error:long_name = "spectral irradiance noise" ;
      		irradiance_error:units = "1" ;
      	byte irradiance_noise(time, scanline, pixel, spectral_channel) ;
      		irradiance_noise:comment = "The irradiance_noise is a measure for the one standard deviation random error of the irradiance measurement; it is expressed in decibel (dB), i.e. 10 times the base-10 logarithmic value of the ratio between the irradiance and the random error." ;
      		irradiance_noise:coordinates = "longitude latitude" ;
      		irradiance_noise:units = "1" ;
      		irradiance_noise:_FillValue = -127b ;
      		irradiance_noise:long_name = "spectral photon irradiance noise, one standard deviation" ;
      	ubyte quality_level(time, scanline, pixel, spectral_channel) ;
      		quality_level:comment = "Overall quality assessment information for each (spectral) pixel" ;
      		quality_level:coordinates = "longitude latitude" ;
      		quality_level:_FillValue = 255UB ;
      		quality_level:long_name = "qualiy level of spectral channel" ;
      		quality_level:max_val = 100UB ;
      		quality_level:min_val = 0UB ;
      		quality_level:units = "mol.m-2.nm-1.s-1" ;
      	ubyte spectral_channel_quality(time, scanline, pixel, spectral_channel) ;
      		spectral_channel_quality:comment = "Quality assessment information for each (spectral) pixel" ;
      		spectral_channel_quality:coordinates = "longitude latitude" ;
      		spectral_channel_quality:_FillValue = 255UB ;
      		spectral_channel_quality:flag_values = 0UB, 1UB, 2UB, 8UB, 16UB, 32UB, 64UB, 128UB ;
      		spectral_channel_quality:flag_masks = 0UB, 1UB, 2UB, 8UB, 16UB, 32UB, 64UB, 128UB ;
      		spectral_channel_quality:flag_meanings = "no_error missing bad_pixel processing_error saturated transient rts underflow" ;
      		spectral_channel_quality:long_name = "spectral channel quality flag" ;
      		spectral_channel_quality:max_val = 254UB ;
      		spectral_channel_quality:min_val = 0UB ;
      		spectral_channel_quality:units = "mol.m-2.nm-1.s-1" ;
      	int time(time) ;
      		time:comment = "Reference time of the measurements. The reference time is set to yyyy-mm-ddT00:00:00 UTC, where yyyy-mm-dd is the day on which the measurements of a particular data granule start." ;
      		time:long_name = "reference start time of measurement" ;
      		time:standard_name = "time" ;
      		time:units = "seconds since 2010-01-01 00:00:00" ;
      } // group OBSERVATIONS

    group: GEODATA {
      variables:
      	float earth_sun_distance(time) ;
      		earth_sun_distance:comment = "1 ua equals 149,597,870,700 meters" ;
      		earth_sun_distance:_FillValue = 9.96921e+36f ;
      		earth_sun_distance:long_name = "distance between the earth and the sun" ;
      		earth_sun_distance:max_val = 1.02f ;
      		earth_sun_distance:min_val = 0.98f ;
      		earth_sun_distance:units = "ua" ;
      } // group GEODATA
    } // group STANDARD_MODE
  } // group BAND4_IRRADIANCE

group: BAND5_IRRADIANCE {

  group: STANDARD_MODE {
    dimensions:
    	time = 1 ;
    	pixel = 308 ;
    	spectral_channel = 497 ;
    	scanline = 1 ;
    	nsettings = 1 ;
    	nbinningregions = 18 ;

    group: OBSERVATIONS {
      variables:
      	int pixel(pixel) ;
      		pixel:comment = "This dimension variable defines the indices across track; index starts at 0" ;
      		pixel:long_name = "across track dimension index" ;
      		pixel:units = "1" ;
      	int spectral_channel(spectral_channel) ;
      		spectral_channel:comment = "This dimension variable defines the indices spectral dimension; index starts at 0" ;
      		spectral_channel:long_name = "wavelength dimension index" ;
      		spectral_channel:units = "1" ;
      	int scanline(scanline) ;
      		scanline:comment = "This dimension variable defines the indices along track; index starts at 0" ;
      		scanline:long_name = "along track dimension index" ;
      		scanline:units = "1" ;
      	int delta_time(time, scanline) ;
      		delta_time:comment = "Time difference with time for each measurement" ;
      		delta_time:_FillValue = -2147483647 ;
      		delta_time:long_name = "offset from the reference start time of measurement" ;
      		delta_time:units = "milliseconds since 2014-08-27 00:00:00" ;
      	ushort detector_column_qualification(time, scanline, spectral_channel) ;
      		detector_column_qualification:comment = "Qualification flag indicating column indicating column type or state" ;
      		detector_column_qualification:_FillValue = 65535US ;
      		detector_column_qualification:flag_values = 0US, 1US, 16US, 32US, 64US, 256US, 512US, 1024US, 2048US ;
      		detector_column_qualification:flag_masks = 0US, 1US, 16US, 98US, 98US, 3840US, 3840US, 3840US, 3840US ;
      		detector_column_qualification:flag_meanings = "no_qualification skipped uvn_odd uvn_prepost uvn_overscan swir_adc0 swir_adc1 swir_adc2 swir_adc3" ;
      		detector_column_qualification:long_name = "Detector column qualification flags" ;
      		detector_column_qualification:max_val = 65534US ;
      		detector_column_qualification:min_val = 0US ;
      		detector_column_qualification:units = "1" ;
      	ushort detector_row_qualification(time, scanline, pixel) ;
      		detector_row_qualification:comment = "Qualification flag indicating row type or state" ;
      		detector_row_qualification:_FillValue = 65535US ;
      		detector_row_qualification:flag_values = 0US, 1US, 2US, 4US, 8US, 16US, 256US, 4096US, 8192US ;
      		detector_row_qualification:flag_masks = 0US, 9US, 2US, 4US, 9US, 16US, 256US, 4096US, 8192US ;
      		detector_row_qualification:flag_meanings = "no_qualification uvn_ror uvn_dump uvn_covered uvn_overscan uvn_higain swir_reference gen_transistion gen_non_illuminated" ;
      		detector_row_qualification:long_name = "Detector row qualification flags" ;
      		detector_row_qualification:max_val = 65534US ;
      		detector_row_qualification:min_val = 0US ;
      		detector_row_qualification:units = "1" ;
      	ushort measurement_quality(time, scanline) ;
      		measurement_quality:flag_values = 0US, 1US, 2US, 16US, 32US, 128US, 256US, 4096US ;
      		measurement_quality:flag_masks = 0US, 1US, 2US, 16US, 32US, 128US, 256US, 4096US ;
      		measurement_quality:flag_meanings = "no_error proc_skipped no_residual saa spacecraft_manoeuvre sub_grp irr_out_of_range sub_group" ;
      		measurement_quality:long_name = "measurement quality flag" ;
      		measurement_quality:max_val = 65534US ;
      		measurement_quality:min_val = 0US ;
      		measurement_quality:units = "1" ;
      		measurement_quality:comment = "Overall quality information for a measurement" ;
      		measurement_quality:coordinates = "longitude latitude" ;
      		measurement_quality:_FillValue = 65535US ;
      	float irradiance(time, scanline, pixel, spectral_channel) ;
      		irradiance:ancilary_vars = "irradiance_noise irradiance_error quality_level spectral_channel_quality" ;
      		irradiance:comment = "Measured spectral irradiance for each spectral pixel" ;
      		irradiance:_FillValue = 9.96921e+36f ;
      		irradiance:long_name = "spectral photon irradiance" ;
      		irradiance:units = "mol.m-2.nm-1.s-1" ;
      	byte irradiance_error(time, scanline, pixel, spectral_channel) ;
      		irradiance_error:comment = "The irradiance_error is a measure for the one standard deviation error of the bias of the irradiance measurement; it is expressed in decibel (dB), i.e. 10 times the base-10 logarithmic value of the ratio between the irradiance and the estimation error." ;
      		irradiance_error:coordinates = "longitude latitude" ;
      		irradiance_error:_FillValue = -127b ;
      		irradiance_error:long_name = "spectral irradiance noise" ;
      		irradiance_error:units = "1" ;
      	byte irradiance_noise(time, scanline, pixel, spectral_channel) ;
      		irradiance_noise:comment = "The irradiance_noise is a measure for the one standard deviation random error of the irradiance measurement; it is expressed in decibel (dB), i.e. 10 times the base-10 logarithmic value of the ratio between the irradiance and the random error." ;
      		irradiance_noise:coordinates = "longitude latitude" ;
      		irradiance_noise:_FillValue = -127b ;
      		irradiance_noise:long_name = "spectral photon irradiance noise, one standard deviation" ;
      		irradiance_noise:units = "1" ;
      	ubyte quality_level(time, scanline, pixel, spectral_channel) ;
      		quality_level:comment = "Overall quality assessment information for each (spectral) pixel" ;
      		quality_level:coordinates = "longitude latitude" ;
      		quality_level:_FillValue = 255UB ;
      		quality_level:long_name = "qualiy level of spectral channel" ;
      		quality_level:max_val = 100UB ;
      		quality_level:min_val = 0UB ;
      		quality_level:units = "mol.m-2.nm-1.s-1" ;
      	ubyte spectral_channel_quality(time, scanline, pixel, spectral_channel) ;
      		spectral_channel_quality:comment = "Quality assessment information for each (spectral) pixel" ;
      		spectral_channel_quality:coordinates = "longitude latitude" ;
      		spectral_channel_quality:_FillValue = 255UB ;
      		spectral_channel_quality:flag_values = 0UB, 1UB, 2UB, 8UB, 16UB, 32UB, 64UB, 128UB ;
      		spectral_channel_quality:flag_masks = 0UB, 1UB, 2UB, 8UB, 16UB, 32UB, 64UB, 128UB ;
      		spectral_channel_quality:flag_meanings = "no_error missing bad_pixel processing_error saturated transient rts underflow" ;
      		spectral_channel_quality:long_name = "spectral channel quality flag" ;
      		spectral_channel_quality:max_val = 254UB ;
      		spectral_channel_quality:min_val = 0UB ;
      		spectral_channel_quality:units = "mol.m-2.nm-1.s-1" ;
      	int time(time) ;
      		time:comment = "Reference time of the measurements. The reference time is set to yyyy-mm-ddT00:00:00 UTC, where yyyy-mm-dd is the day on which the measurements of a particular data granule start." ;
      		time:long_name = "reference start time of measurement" ;
      		time:standard_name = "time" ;
      		time:units = "seconds since 2010-01-01 00:00:00" ;
      } // group OBSERVATIONS

    group: GEODATA {
      variables:
      	float earth_sun_distance(time) ;
      		earth_sun_distance:comment = "1 ua equals 149,597,870,700 meters" ;
      		earth_sun_distance:_FillValue = 9.96921e+36f ;
      		earth_sun_distance:long_name = "distance between the earth and the sun" ;
      		earth_sun_distance:max_val = 1.02f ;
      		earth_sun_distance:min_val = 0.98f ;
      		earth_sun_distance:units = "ua" ;
      } // group GEODATA
    } // group STANDARD_MODE
  } // group BAND5_IRRADIANCE

group: BAND6_IRRADIANCE {

  group: STANDARD_MODE {
    dimensions:
    	time = 1 ;
    	pixel = 448 ;
    	spectral_channel = 497 ;
    	scanline = 1 ;
    	nsettings = 1 ;
    	nbinningregions = 18 ;

    group: OBSERVATIONS {
      variables:
      	int pixel(pixel) ;
      		pixel:comment = "This dimension variable defines the indices across track; index starts at 0" ;
      		pixel:long_name = "across track dimension index" ;
      		pixel:units = "1" ;
      	int spectral_channel(spectral_channel) ;
      		spectral_channel:comment = "This dimension variable defines the indices spectral dimension; index starts at 0" ;
      		spectral_channel:long_name = "wavelength dimension index" ;
      		spectral_channel:units = "1" ;
      	int scanline(scanline) ;
      		scanline:comment = "This dimension variable defines the indices along track; index starts at 0" ;
      		scanline:long_name = "along track dimension index" ;
      		scanline:units = "1" ;
      	int delta_time(time, scanline) ;
      		delta_time:comment = "Time difference with time for each measurement" ;
      		delta_time:_FillValue = -2147483647 ;
      		delta_time:long_name = "offset from the reference start time of measurement" ;
      		delta_time:units = "milliseconds since 2014-08-27 00:00:00" ;
      	ushort detector_column_qualification(time, scanline, spectral_channel) ;
      		detector_column_qualification:comment = "Qualification flag indicating column indicating column type or state" ;
      		detector_column_qualification:_FillValue = 65535US ;
      		detector_column_qualification:flag_values = 0US, 1US, 16US, 32US, 64US, 256US, 512US, 1024US, 2048US ;
      		detector_column_qualification:flag_masks = 0US, 1US, 16US, 98US, 98US, 3840US, 3840US, 3840US, 3840US ;
      		detector_column_qualification:flag_meanings = "no_qualification skipped uvn_odd uvn_prepost uvn_overscan swir_adc0 swir_adc1 swir_adc2 swir_adc3" ;
      		detector_column_qualification:long_name = "Detector column qualification flags" ;
      		detector_column_qualification:max_val = 65534US ;
      		detector_column_qualification:min_val = 0US ;
      		detector_column_qualification:units = "1" ;
      	ushort detector_row_qualification(time, scanline, pixel) ;
      		detector_row_qualification:comment = "Qualification flag indicating row type or state" ;
      		detector_row_qualification:_FillValue = 65535US ;
      		detector_row_qualification:flag_values = 0US, 1US, 2US, 4US, 8US, 16US, 256US, 4096US, 8192US ;
      		detector_row_qualification:flag_masks = 0US, 9US, 2US, 4US, 9US, 16US, 256US, 4096US, 8192US ;
      		detector_row_qualification:flag_meanings = "no_qualification uvn_ror uvn_dump uvn_covered uvn_overscan uvn_higain swir_reference gen_transistion gen_non_illuminated" ;
      		detector_row_qualification:long_name = "Detector row qualification flags" ;
      		detector_row_qualification:max_val = 65534US ;
      		detector_row_qualification:min_val = 0US ;
      		detector_row_qualification:units = "1" ;
      	ushort measurement_quality(time, scanline) ;
      		measurement_quality:flag_values = 0US, 1US, 2US, 16US, 32US, 128US, 256US, 4096US ;
      		measurement_quality:flag_masks = 0US, 1US, 2US, 16US, 32US, 128US, 256US, 4096US ;
      		measurement_quality:flag_meanings = "no_error proc_skipped no_residual saa spacecraft_manoeuvre sub_grp irr_out_of_range sub_group" ;
      		measurement_quality:long_name = "measurement quality flag" ;
      		measurement_quality:max_val = 65534US ;
      		measurement_quality:min_val = 0US ;
      		measurement_quality:units = "1" ;
      		measurement_quality:comment = "Overall quality information for a measurement" ;
      		measurement_quality:coordinates = "longitude latitude" ;
      		measurement_quality:_FillValue = 65535US ;
      	float irradiance(time, scanline, pixel, spectral_channel) ;
      		irradiance:ancilary_vars = "irradiance_noise irradiance_error quality_level spectral_channel_quality" ;
      		irradiance:comment = "Measured spectral irradiance for each spectral pixel" ;
      		irradiance:_FillValue = 9.96921e+36f ;
      		irradiance:long_name = "spectral photon irradiance" ;
      		irradiance:units = "mol.m-2.nm-1.s-1" ;
      	byte irradiance_error(time, scanline, pixel, spectral_channel) ;
      		irradiance_error:comment = "The irradiance_error is a measure for the one standard deviation error of the bias of the irradiance measurement; it is expressed in decibel (dB), i.e. 10 times the base-10 logarithmic value of the ratio between the irradiance and the estimation error." ;
      		irradiance_error:coordinates = "longitude latitude" ;
      		irradiance_error:_FillValue = -127b ;
      		irradiance_error:long_name = "spectral irradiance noise" ;
      		irradiance_error:units = "1" ;
      	byte irradiance_noise(time, scanline, pixel, spectral_channel) ;
      		irradiance_noise:comment = "The irradiance_noise is a measure for the one standard deviation random error of the irradiance measurement; it is expressed in decibel (dB), i.e. 10 times the base-10 logarithmic value of the ratio between the irradiance and the random error." ;
      		irradiance_noise:coordinates = "longitude latitude" ;
      		irradiance_noise:units = "1" ;
      		irradiance_noise:_FillValue = -127b ;
      		irradiance_noise:long_name = "spectral photon irradiance noise, one standard deviation" ;
      	ubyte quality_level(time, scanline, pixel, spectral_channel) ;
      		quality_level:comment = "Overall quality assessment information for each (spectral) pixel" ;
      		quality_level:coordinates = "longitude latitude" ;
      		quality_level:_FillValue = 255UB ;
      		quality_level:long_name = "qualiy level of spectral channel" ;
      		quality_level:max_val = 100UB ;
      		quality_level:min_val = 0UB ;
      		quality_level:units = "mol.m-2.nm-1.s-1" ;
      	ubyte spectral_channel_quality(time, scanline, pixel, spectral_channel) ;
      		spectral_channel_quality:comment = "Quality assessment information for each (spectral) pixel" ;
      		spectral_channel_quality:coordinates = "longitude latitude" ;
      		spectral_channel_quality:_FillValue = 255UB ;
      		spectral_channel_quality:flag_values = 0UB, 1UB, 2UB, 8UB, 16UB, 32UB, 64UB, 128UB ;
      		spectral_channel_quality:max_val = 254UB ;
      		spectral_channel_quality:flag_masks = 0UB, 1UB, 2UB, 8UB, 16UB, 32UB, 64UB, 128UB ;
      		spectral_channel_quality:flag_meanings = "no_error missing bad_pixel processing_error saturated transient rts underflow" ;
      		spectral_channel_quality:long_name = "spectral channel quality flag" ;
      		spectral_channel_quality:min_val = 0UB ;
      		spectral_channel_quality:units = "mol.m-2.nm-1.s-1" ;
      	int time(time) ;
      		time:comment = "Reference time of the measurements. The reference time is set to yyyy-mm-ddT00:00:00 UTC, where yyyy-mm-dd is the day on which the measurements of a particular data granule start." ;
      		time:long_name = "reference start time of measurement" ;
      		time:standard_name = "time" ;
      		time:units = "seconds since 2010-01-01 00:00:00" ;
      } // group OBSERVATIONS

    group: GEODATA {
      variables:
      	float earth_sun_distance(time) ;
      		earth_sun_distance:comment = "1 ua equals 149,597,870,700 meters" ;
      		earth_sun_distance:_FillValue = 9.96921e+36f ;
      		earth_sun_distance:long_name = "distance between the earth and the sun" ;
      		earth_sun_distance:max_val = 1.02f ;
      		earth_sun_distance:min_val = 0.98f ;
      		earth_sun_distance:units = "ua" ;
      } // group GEODATA
    } // group STANDARD_MODE
  } // group BAND6_IRRADIANCE
}
