// Provided by Jim Biard, jbiard@cicsnc.org
//
// This example is an attempt to produce a NOAA Level 1b file using netCDF. The
// file contains everything needed to reproduce the original CCSDS downlink
// data packets (Level 1a). It is a "superuser" data set, in that the intended
// audience is reprocessors. All measurements have been demultiplexed and
// stored as separate variables according to their kind.
//
//
netcdf CVIRS_npp_d20160606_t0707464_e0713278_b23876_c20160606220333548229_ncdc_ops {
dimensions:
	scans = UNLIMITED ; // (192 currently)
	granules = UNLIMITED ; // (4 currently)

// global attributes:
		string :acknowledgment = "This project was supported by the NOAA Climate Data Record (CDR) Program for satellites." ;
		string :cdm_data_type = "SWATH" ;
		string :Conventions = "CF-1.5" ;
		string :creator_url = "http://www.ncdc.noaa.gov" ;
		string :geospatial_lat_units = "degrees_east" ;
		string :geospatial_lon_units = "degrees_north" ;
		string :history = "Initial release" ;
		string :institution = "DOC/NOAA/NESDIS/NCDC > National Climatic Data Center, NESDIS, NOAA, U.S. Department of Commerce" ;
		string :keywords = "EARTH SCIENCE > SPECTRAL/ENGINEERING > VISIBLE WAVELENGTHS > SENSOR COUNTS, EARTH SCIENCE > SPECTRAL/ENGINEERING > PLATFORM CHARACTERISTICS > AIRSPEED/GROUND SPEED, EARTH SCIENCE > SPECTRAL/ENGINEERING > PLATFORM CHARACTERISTICS > ATTITUDE CHARACTERISTICS, EARTH SCIENCE > SPECTRAL/ENGINEERING > PLATFORM CHARACTERISTICS > DATA SYNCHRONIZATION TIME, EARTH SCIENCE > SPECTRAL/ENGINEERING > PLATFORM CHARACTERISTICS > ORBITAL CHARACTERISTICS, EARTH SCIENCE > SPECTRAL/ENGINEERING > PLATFORM CHARACTERISTICS > VIEWING GEOMETRY, EARTH SCIENCE > SPECTRAL/ENGINEERING > SENSOR CHARACTERISTICS > ELECTRICAL PROPERTIES, EARTH SCIENCE > SPECTRAL/ENGINEERING > SENSOR CHARACTERISTICS > PHASE AND AMPLITUDE, EARTH SCIENCE > SPECTRAL/ENGINEERING > SENSOR CHARACTERISTICS > THERMAL PROPERTIES, EARTH SCIENCE > SPECTRAL/ENGINEERING > SENSOR CHARACTERISTICS > TOTAL TEMPERATURE, EARTH SCIENCE > SPECTRAL/ENGINEERING > SENSOR CHARACTERISTICS > VIEWING GEOMETRY" ;
		string :keywords_vocabulary = "NASA Global Change Master Directory (GCMD) Science Keywords, Version 7.0" ;
		string :license = "No constraints on data access or use." ;
		string :Metadata_Conventions = "CF-1.6, Unidata Dataset Discovery v1.0, Suomi NPP CDFCB-X, Suomi NPP MDFCB" ;
		string :Metadata_Link = "gov.noaa.ncdc:C00836" ;
		string :naming_authority = "DOC/NOAA/NESDIS/NCDC > National Climatic Data Center, NESDIS, NOAA, U.S. Department of Commerce" ;
		string :processing_level = "NOAA Level 1b" ;
		string :publisher_name = "DOC/NOAA/NESDIS/NCDC > National Climatic Data Center, NESDIS, NOAA, U.S. Department of Commerce" ;
		string :publisher_url = "http://www.ncdc.noaa.gov" ;
		string :standard_name_vocabulary = "CF Standard Name Table (v22, 12 February 2013)" ;
		string :summary = "The Suomi NPP Climate Raw Data Record (C-RDR) is an intermediate processing level (level 1b) between a Raw Data Record and a Sensor Data Record. The C-RDR is intended to simplify access to the raw data for the purpose of reprocessing using calibration and geolocation methods. This C-RDR has raw Visible Infrared Imager Radiometer Suite (VIIRS) measurements collected into time series variables, accompanied by the coefficients and tables needed to convert them to science units and calibrate them. The measurements, processing coefficients, and LUTs are stored as variables organized into netCDF-4 groups. The netCDF-4 groups are Engineering_Data, Image_375m, Image_750m_DualGain, Image_750m_SingleGain, Image_DayNight, Quality_Measures, and Spacecraft_Diary. Where applicable, metadata in this file follows the Climate and Forecast (CF) Conventions and Attribute Convention for Dataset Discovery (ACDD). Metadata attributes from the native Suomi NPP RDR and SDR file types are also included. These files have been compared with those generated using JPSS Application Development Library (ADL) applications." ;
		string :title = "Suomi-NPP VIIRS C-RDR (Draft)" ;
		string :Processing_Software_ID = "TBD" ;
		string :Processing_Software_Version = "TBD" ;
		string :references = "VIIRS C-RDR Product Specification (CDRP-EXT-0247), JPSS Common Data Format Control Book - External (CDFCB-X) (474-00001), NPP Mission Data Format Control Book (MDFCB) (GSFC 429-05-02-42)" ;
		string :missing_value_meanings = "ScaleOutOfBounds ValueDoesNotExist EllipsoidIntersectionFailed CannotCalculate OnGroundPixelTrim OnBoardPixelTrim Missing NotApplicable" ;
		string :missing_values_8bit_signed = "120 121 122 123 124 125 126 127" ;
		string :missing_values_8bit_unsigned = "248 249 250 251 252 253 254 255" ;
		string :missing_values_16bit_signed = "-992 -993 -994 -995 -996 -997 -998 -999" ;
		string :missing_values_16bit_unsigned = "65528 65529 65530 65531 65532 65533 65534 65535" ;
		string :missing_values_32bit_signed = "-992 -993 -994 -995 -996 -997 -998 -999" ;
		string :missing_values_32bit_unsigned = "4294967288 4294967289 4294967290 4294967291 4294967292 4294967293 4294967294 4294967295" ;
		string :missing_values_64bit_signed = "-992 -993 -994 -995 -996 -997 -998 -999" ;
		string :missing_values_64bit_unsigned = "18446744073709551608 18446744073709551609 18446744073709551610 18446744073709551611 18446744073709551612 18446744073709551613 18446744073709551614 18446744073709551615" ;
		string :missing_values_32bit_float = "-999.2 -999.3 -999.4 -999.5 -999.6 -999.7 -999.8 -999.9" ;
		string :missing_values_64bit_float = "-999.2 -999.3 -999.4 -999.5 -999.6 -999.7 -999.8 -999.9" ;
		string :date_created = "2016-06-06T22:03:33.548229Z" ;
		string :date_issued = "2016-06-06T22:03:33.548229Z" ;
		string :date_modified = "2016-06-06T22:03:33.548229Z" ;
		:geospatial_lat_max = -51.6182010959577 ;
		:geospatial_lat_min = -77.9912603523064 ;
		:geospatial_lon_max = -57.9768171062649 ;
		:geospatial_lon_min = -151.566223449375 ;
		string :id = "CVIRS_npp_d20160606_t0707464_e0713278_b23876_c20160606220333548229_ncdc_ops.nc" ;
		string :project = "NPP" ;
		string :time_coverage_end = "2016-06-06T07:13:27.850000Z" ;
		string :time_coverage_start = "2016-06-06T07:07:46.450000Z" ;
		string :Ascending_Descending_Indicator = "1", "1", "1", "1" ;
		:Beginning_Orbit_Numbers = 23876, 23876, 23876, 23876 ;
		:Beginning_Time_IET = 1.84388810245e+15 ;
		string :Day_Night_Flag = "Night", "Night", "Night", "Night" ;
		:Ending_Orbit_Number = 23876 ;
		:Ending_Time_IET = 1.84388844385e+15 ;
		:GRing_Latitudes = -51.6182010959577, -53.5907977929865, -55.5748470394461, -57.2972287000934, -59.0976507177469, -60.6244689092769, -62.1753814427987, -63.4319898536618, -64.6438781283422, -76.0843399427066, -77.9912603523064, -75.6680460472547, -73.373042905582, -71.0608666756226, -68.6933960365745, -66.3312223692378, -63.9279752777636, -61.538434096537, -59.1144885037355, -57.9344442840345, -51.6182010959577 ;
		:GRing_Longitudes = -121.687139610264, -124.246982861944, -127.20717941289, -130.178410050814, -133.795236336388, -137.429304109931, -141.841910157803, -146.258135279347, -151.566223449375, -124.843434367837, -57.9768171062649, -62.4180287378294, -65.363657108712, -67.4708321566642, -69.0495060554353, -70.2118730377681, -71.1059770083863, -71.7621760535086, -72.265872052918, -99.5318997887377, -121.687139610264 ;
		string :Input_RDR_Granule_IDs = "NPP001458688684", "NPP001458689538", "NPP001458690391", "NPP001458691245" ;
		string :Input_RDR_Granule_Versions = "A1", "A1", "A1", "A1" ;
		string :Input_Support_File_IDs = "off_Planet-Eph-ANC_Static_JPL_000f_20000101_200001010000Z_20000101000000Z_ee00000000000000Z_np", "CMNGEO-PARAM-LUT_npp_20020101010000Z_20020101010000Z_ee00000000000000Z_PS-1-D-NPP-1-PE-_devl_dev_all-_all", "VIIRS-SDR-GEO-DNB-PARAM-LUT_npp_20020101010000Z_20020101010000Z_ee00000000000000Z_PS-1-D-NPP-5-PE-_devl_dev_all-_all", "VIIRS-SDR-GEO-IMG-PARAM-LUT_npp_20020101010000Z_20020101010000Z_ee00000000000000Z_PS-1-D-NPP-5-PE-_devl_dev_all-_all", "VIIRS-SDR-GEO-MOD-PARAM-LUT_npp_20020101010000Z_20020101010000Z_ee00000000000000Z_PS-1-D-NPP-5-PE-_devl_dev_all-_all", "VIIRS-SDR-QA-LUT_npp_20020101010000Z_20020101010000Z_ee00000000000000Z_1_devl_dev_all-_all" ;
		string :Instrument = "VIIRS" ;
		string :Instrument_Flight_Software_Version = "23" ;
		string :LEOA_Flags = "Off", "Off", "Off", "Off" ;
		:Nadir_Latitude_Max = -57.9849801538946 ;
		:Nadir_Latitude_Min = -76.0408054605633 ;
		:Nadir_Longitude_Max = -99.5699970661005 ;
		:Nadir_Longitude_Min = -124.723563758053 ;
		string :NPP_Processing_Domain_ID = "ops" ;
		:Number_Of_Scans = 192 ;
		string :Operational_Mode = "NPP Unknown, VIIRS Operational", "NPP Unknown, VIIRS Operational", "NPP Unknown, VIIRS Operational", "NPP Unknown, VIIRS Operational" ;
		:Percent_Erroneous_Data = 0. ;
		:Percent_Missing_Data = 0. ;
		:Percent_Not_Applicable_Data = 0. ;
		string :Platform = "NPP" ;
		string :Quality_Summary_Names = "BadChecksum", "DiscardedPackets", "MissingPackets", "PoorQualityScans" ;
		:Quality_Summary_Values = 0., 0., 45120., 0. ;
		:Satellite_Local_Azimuth_Angle_Max = 153.68756236958 ;
		:Satellite_Local_Azimuth_Angle_Min = -158.191048226664 ;
		:Satellite_Local_Zenith_Angle_Max = 70.5977345937329 ;
		:Satellite_Local_Zenith_Angle_Min = 0.0442650909208163 ;
		:Solar_Azimuth_Angle_Max = 179.566811620914 ;
		:Solar_Azimuth_Angle_Min = -176.927073497122 ;
		:Solar_Zenith_Angle_Max = 149.011310656009 ;
		:Solar_Zenith_Angle_Min = 119.9374159056 ;
		string :Spacecraft_Maneuver = "Unknown", "Unknown", "Unknown", "Unknown" ;

group: Engineering_Data {
  dimensions:
  	hrdt_samples = 16 ;
  	mirror_sides = 2 ;
  	encoder_samples = 1290 ;
  	detectors_375m = 32 ;
  	sdsm_detectors_750m = 8 ;
  	sdsm_samples = 5 ;
  	bb_thermistors = 6 ;
  	detectors_750m = 16 ;
  	events = 64 ;
  	event_bytes = 18 ;
  variables:
  	int scans_per_granule(granules) ;
  		scans_per_granule:_FillValue = -998 ;
  		scans_per_granule:valid_min = -2147483648 ;
  		scans_per_granule:valid_max = 2147483647 ;
  		scans_per_granule:missing_value = -992, -993, -994, -995, -996, -997, -998, -999 ;
  		string scans_per_granule:long_name = "Number of scans for each granule" ;
  	int starting_scan_per_granule(granules) ;
  		starting_scan_per_granule:_FillValue = -998 ;
  		starting_scan_per_granule:valid_min = -2147483648 ;
  		starting_scan_per_granule:valid_max = 2147483647 ;
  		starting_scan_per_granule:missing_value = -992, -993, -994, -995, -996, -997, -998, -999 ;
  		string starting_scan_per_granule:long_name = "Index of the scan that starts each granule" ;
  	double start_of_scan_time(scans) ;
  		start_of_scan_time:_FillValue = -999.8 ;
  		start_of_scan_time:valid_min = 1.48323e+15 ;
  		start_of_scan_time:valid_max = 2.27215e+15 ;
  		start_of_scan_time:missing_value = -999.2, -999.3, -999.4, -999.5, -999.6, -999.7, -999.8, -999.9 ;
  		string start_of_scan_time:units = "microseconds since 1958/01/01 00:00:00" ;
  		string start_of_scan_time:long_name = "Scan Start Time" ;
  		string start_of_scan_time:source = "APID826:SecondaryHeader.StartOfScan" ;
  		string start_of_scan_time:standard_name = "time" ;
  	uint s_cp_seq_cnt(scans) ;
  		s_cp_seq_cnt:_FillValue = 4294967294U ;
  		s_cp_seq_cnt:valid_min = 0U ;
  		s_cp_seq_cnt:valid_max = 4294967295U ;
  		s_cp_seq_cnt:missing_value = 4294967288U, 0U, 4294967289U, 0U, 4294967290U, 0U, 4294967291U, 0U ;
  		string s_cp_seq_cnt:coordinates = "start_of_scan_time" ;
  		string s_cp_seq_cnt:long_name = "Total Packet Count" ;
  		string s_cp_seq_cnt:source = "APID826:S_CP_SEQ_CNT" ;
  	double s_cp_pkt_time(scans) ;
  		s_cp_pkt_time:_FillValue = -999.8 ;
  		s_cp_pkt_time:valid_min = 1.48323e+15 ;
  		s_cp_pkt_time:valid_max = 2.27215e+15 ;
  		s_cp_pkt_time:missing_value = -999.2, -999.3, -999.4, -999.5, -999.6, -999.7, -999.8, -999.9 ;
  		string s_cp_pkt_time:coordinates = "start_of_scan_time" ;
  		string s_cp_pkt_time:units = "microseconds since 1958/01/01 00:00:00" ;
  		string s_cp_pkt_time:long_name = "Packet Time" ;
  		string s_cp_pkt_time:source = "APID826:(S_CP_PKT_TIME_DAY, S_CP_PKT_TIME_MILLISEC, S_CP_PKT_TIME_MICROSEC)" ;
  		string s_cp_pkt_time:standard_name = "time" ;
  	ubyte c_cp_format_ver(scans) ;
  		c_cp_format_ver:_FillValue = 254UB ;
  		c_cp_format_ver:valid_min = 1UB ;
  		c_cp_format_ver:valid_max = 248UB ;
  		c_cp_format_ver:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string c_cp_format_ver:coordinates = "start_of_scan_time" ;
  		string c_cp_format_ver:long_name = "Telemetry Format Version" ;
  		string c_cp_format_ver:source = "APID826:C_CP_FORMAT_VER" ;
  	ubyte c_cp_instr_num(scans) ;
  		c_cp_instr_num:_FillValue = 254UB ;
  		c_cp_instr_num:valid_min = 1UB ;
  		c_cp_instr_num:valid_max = 248UB ;
  		c_cp_instr_num:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string c_cp_instr_num:coordinates = "start_of_scan_time" ;
  		string c_cp_instr_num:long_name = "Instrument ID" ;
  		string c_cp_instr_num:source = "APID826:C_CP_INSTR_NUM" ;
  	ushort c_cp_fsw_version(scans) ;
  		c_cp_fsw_version:_FillValue = 65534US ;
  		c_cp_fsw_version:valid_min = 12289US ;
  		c_cp_fsw_version:valid_max = 32767US ;
  		c_cp_fsw_version:missing_value = 65528US, 65529US, 65530US, 65531US, 65532US, 65533US, 65534US, 65535US ;
  		string c_cp_fsw_version:coordinates = "start_of_scan_time" ;
  		string c_cp_fsw_version:long_name = "Flight Hardware and Software Version" ;
  		string c_cp_fsw_version:source = "APID826:C_CP_FSW_VERSION" ;
  	double s_cp_end_scan_time(scans) ;
  		s_cp_end_scan_time:_FillValue = -999.8 ;
  		s_cp_end_scan_time:valid_min = 1.48323e+15 ;
  		s_cp_end_scan_time:valid_max = 2.27215e+15 ;
  		s_cp_end_scan_time:missing_value = -999.2, -999.3, -999.4, -999.5, -999.6, -999.7, -999.8, -999.9 ;
  		string s_cp_end_scan_time:coordinates = "start_of_scan_time" ;
  		string s_cp_end_scan_time:units = "microseconds since 1958/01/01 00:00:00" ;
  		string s_cp_end_scan_time:long_name = "Scan End Time" ;
  		string s_cp_end_scan_time:source = "APID826:(S_CP_END_SCAN_DAY, S_CP_END_SCAN_MILLISEC, S_CP_END_SCAN_MICROSEC)" ;
  		string s_cp_end_scan_time:standard_name = "time" ;
  	uint s_cp_scan_num(scans) ;
  		s_cp_scan_num:_FillValue = 4294967294U ;
  		s_cp_scan_num:valid_min = 0U ;
  		s_cp_scan_num:valid_max = 4294967295U ;
  		s_cp_scan_num:missing_value = 4294967288U, 0U, 4294967289U, 0U, 4294967290U, 0U, 4294967291U, 0U ;
  		string s_cp_scan_num:coordinates = "start_of_scan_time" ;
  		string s_cp_scan_num:long_name = "Scan Number" ;
  		string s_cp_scan_num:source = "APID826:S_CP_SCAN_NUM" ;
  	ubyte s_cp_sensor_mode(scans) ;
  		s_cp_sensor_mode:_FillValue = 254UB ;
  		s_cp_sensor_mode:valid_min = 0UB ;
  		s_cp_sensor_mode:valid_max = 7UB ;
  		s_cp_sensor_mode:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string s_cp_sensor_mode:coordinates = "start_of_scan_time" ;
  		string s_cp_sensor_mode:long_name = "Sensor Mode" ;
  		string s_cp_sensor_mode:source = "APID826:S_CP_SENSOR_MODE" ;
  	ubyte s_cp_servo_locked(scans) ;
  		s_cp_servo_locked:_FillValue = 254UB ;
  		s_cp_servo_locked:valid_min = 0UB ;
  		s_cp_servo_locked:valid_max = 1UB ;
  		s_cp_servo_locked:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string s_cp_servo_locked:coordinates = "start_of_scan_time" ;
  		string s_cp_servo_locked:long_name = "Servo Locked" ;
  		string s_cp_servo_locked:source = "APID826:S_CP_SERVO_LOCKED" ;
  	ubyte s_cp_ham_side(scans) ;
  		s_cp_ham_side:_FillValue = 254UB ;
  		s_cp_ham_side:valid_min = 0UB ;
  		s_cp_ham_side:valid_max = 1UB ;
  		s_cp_ham_side:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string s_cp_ham_side:coordinates = "start_of_scan_time" ;
  		string s_cp_ham_side:long_name = "Half Angle Mirror Side" ;
  		string s_cp_ham_side:source = "APID826:S_CP_HAM_SIDE" ;
  	ubyte s_cp_sdsm_active(scans) ;
  		s_cp_sdsm_active:_FillValue = 254UB ;
  		s_cp_sdsm_active:valid_min = 0UB ;
  		s_cp_sdsm_active:valid_max = 1UB ;
  		s_cp_sdsm_active:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string s_cp_sdsm_active:coordinates = "start_of_scan_time" ;
  		string s_cp_sdsm_active:long_name = "SDSM Active" ;
  		string s_cp_sdsm_active:source = "APID826:S_CP_SDSM_ACTIVE" ;
  	ubyte s_cp_fpa_cal_data_gain(scans) ;
  		s_cp_fpa_cal_data_gain:_FillValue = 254UB ;
  		s_cp_fpa_cal_data_gain:valid_min = 0UB ;
  		s_cp_fpa_cal_data_gain:valid_max = 1UB ;
  		s_cp_fpa_cal_data_gain:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string s_cp_fpa_cal_data_gain:coordinates = "start_of_scan_time" ;
  		string s_cp_fpa_cal_data_gain:long_name = "FPA Calibration Data Gain" ;
  		string s_cp_fpa_cal_data_gain:source = "APID826:S_CP_FPA_CAL_DATA_GAIN" ;
  	ubyte s_cp_self_test_data(scans) ;
  		s_cp_self_test_data:_FillValue = 254UB ;
  		s_cp_self_test_data:valid_min = 0UB ;
  		s_cp_self_test_data:valid_max = 15UB ;
  		s_cp_self_test_data:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string s_cp_self_test_data:coordinates = "start_of_scan_time" ;
  		string s_cp_self_test_data:long_name = "Self-test Data Pattern" ;
  		string s_cp_self_test_data:source = "APID826:S_CP_SELF_TEST_DATA" ;
  	ubyte es_se_a_teleham_scansync(scans) ;
  		es_se_a_teleham_scansync:_FillValue = 254UB ;
  		es_se_a_teleham_scansync:valid_min = 0UB ;
  		es_se_a_teleham_scansync:valid_max = 1UB ;
  		es_se_a_teleham_scansync:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string es_se_a_teleham_scansync:coordinates = "start_of_scan_time" ;
  		string es_se_a_teleham_scansync:long_name = "SCE-A Telescope/Half-Angle Mirror Scan Sync" ;
  		string es_se_a_teleham_scansync:source = "APID826:ES_SE_A_TELEHAM_SCANSYN" ;
  	ubyte es_se_b_teleham_scansync(scans) ;
  		es_se_b_teleham_scansync:_FillValue = 254UB ;
  		es_se_b_teleham_scansync:valid_min = 0UB ;
  		es_se_b_teleham_scansync:valid_max = 1UB ;
  		es_se_b_teleham_scansync:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string es_se_b_teleham_scansync:coordinates = "start_of_scan_time" ;
  		string es_se_b_teleham_scansync:long_name = "SCE-B Telescope/Half-Angle Mirror Scan Sync" ;
  		string es_se_b_teleham_scansync:source = "APID826:ES_SE_B_TELEHAM_SCANSYN" ;
  	ubyte es_sd_sdsm_mtr_step_cnt(scans) ;
  		es_sd_sdsm_mtr_step_cnt:_FillValue = 254UB ;
  		es_sd_sdsm_mtr_step_cnt:valid_min = 0UB ;
  		es_sd_sdsm_mtr_step_cnt:valid_max = 127UB ;
  		es_sd_sdsm_mtr_step_cnt:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string es_sd_sdsm_mtr_step_cnt:coordinates = "start_of_scan_time" ;
  		string es_sd_sdsm_mtr_step_cnt:long_name = "SDSM Motor Absolute Step Count" ;
  		string es_sd_sdsm_mtr_step_cnt:source = "APID826:ES_SD_SDSM_MTR_STEP_CNT" ;
  	ubyte c_dp_reg_tbl_rev(scans) ;
  		c_dp_reg_tbl_rev:_FillValue = 254UB ;
  		c_dp_reg_tbl_rev:valid_min = 0UB ;
  		c_dp_reg_tbl_rev:valid_max = 248UB ;
  		c_dp_reg_tbl_rev:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string c_dp_reg_tbl_rev:coordinates = "start_of_scan_time" ;
  		string c_dp_reg_tbl_rev:long_name = "DPP Register Table Revision" ;
  		string c_dp_reg_tbl_rev:source = "APID826:C_DP_REG_TBL_REV" ;
  	ubyte c_dp_state_tran_tbl_rev(scans) ;
  		c_dp_state_tran_tbl_rev:_FillValue = 254UB ;
  		c_dp_state_tran_tbl_rev:valid_min = 0UB ;
  		c_dp_state_tran_tbl_rev:valid_max = 248UB ;
  		c_dp_state_tran_tbl_rev:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string c_dp_state_tran_tbl_rev:coordinates = "start_of_scan_time" ;
  		string c_dp_state_tran_tbl_rev:long_name = "DPP State Transition Table Revision" ;
  		string c_dp_state_tran_tbl_rev:source = "APID826:C_DP_STATE_TRAN_TBL_REV" ;
  	ubyte c_dp_band_proc_tbl_rev(scans) ;
  		c_dp_band_proc_tbl_rev:_FillValue = 254UB ;
  		c_dp_band_proc_tbl_rev:valid_min = 0UB ;
  		c_dp_band_proc_tbl_rev:valid_max = 248UB ;
  		c_dp_band_proc_tbl_rev:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string c_dp_band_proc_tbl_rev:coordinates = "start_of_scan_time" ;
  		string c_dp_band_proc_tbl_rev:long_name = "DPP Band Processing Table Revision" ;
  		string c_dp_band_proc_tbl_rev:source = "APID826:C_DP_BAND_PROC_TBL_REV" ;
  	ubyte c_dp_heat_ctrl_tbl_rev(scans) ;
  		c_dp_heat_ctrl_tbl_rev:_FillValue = 254UB ;
  		c_dp_heat_ctrl_tbl_rev:valid_min = 0UB ;
  		c_dp_heat_ctrl_tbl_rev:valid_max = 248UB ;
  		c_dp_heat_ctrl_tbl_rev:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string c_dp_heat_ctrl_tbl_rev:coordinates = "start_of_scan_time" ;
  		string c_dp_heat_ctrl_tbl_rev:long_name = "PWM Heater Control Table Revision" ;
  		string c_dp_heat_ctrl_tbl_rev:source = "APID826:C_DP_HEAT_CTRL_TBL_REV" ;
  	ubyte c_dp_macro_cmd_tbl_rev(scans) ;
  		c_dp_macro_cmd_tbl_rev:_FillValue = 254UB ;
  		c_dp_macro_cmd_tbl_rev:valid_min = 0UB ;
  		c_dp_macro_cmd_tbl_rev:valid_max = 248UB ;
  		c_dp_macro_cmd_tbl_rev:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string c_dp_macro_cmd_tbl_rev:coordinates = "start_of_scan_time" ;
  		string c_dp_macro_cmd_tbl_rev:long_name = "Macro Command Table Revision" ;
  		string c_dp_macro_cmd_tbl_rev:source = "APID826:C_DP_MACRO_CMD_TBL_REV" ;
  	ubyte c_dp_crit_tele_tbl_rev(scans) ;
  		c_dp_crit_tele_tbl_rev:_FillValue = 254UB ;
  		c_dp_crit_tele_tbl_rev:valid_min = 0UB ;
  		c_dp_crit_tele_tbl_rev:valid_max = 248UB ;
  		c_dp_crit_tele_tbl_rev:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string c_dp_crit_tele_tbl_rev:coordinates = "start_of_scan_time" ;
  		string c_dp_crit_tele_tbl_rev:long_name = "Critical Telemetry Table Revision" ;
  		string c_dp_crit_tele_tbl_rev:source = "APID826:C_DP_CRIT_TELE_TBL_REV" ;
  	ushort c_dp_stor_cmd_tbl_rev(scans) ;
  		c_dp_stor_cmd_tbl_rev:_FillValue = 65534US ;
  		c_dp_stor_cmd_tbl_rev:valid_min = 0US ;
  		c_dp_stor_cmd_tbl_rev:valid_max = 65528US ;
  		c_dp_stor_cmd_tbl_rev:missing_value = 65528US, 65529US, 65530US, 65531US, 65532US, 65533US, 65534US, 65535US ;
  		string c_dp_stor_cmd_tbl_rev:coordinates = "start_of_scan_time" ;
  		string c_dp_stor_cmd_tbl_rev:long_name = "Stored Command Table Revision" ;
  		string c_dp_stor_cmd_tbl_rev:source = "APID826:C_DP_STOR_CMD_TBL_REV" ;
  	ubyte ec_dp_dn_m_l_gain_pkt(scans) ;
  		ec_dp_dn_m_l_gain_pkt:_FillValue = 254UB ;
  		ec_dp_dn_m_l_gain_pkt:valid_min = 0UB ;
  		ec_dp_dn_m_l_gain_pkt:valid_max = 1UB ;
  		ec_dp_dn_m_l_gain_pkt:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string ec_dp_dn_m_l_gain_pkt:coordinates = "start_of_scan_time" ;
  		string ec_dp_dn_m_l_gain_pkt:long_name = "Send Day/Night Band Low and Middle Gain Stage Packets" ;
  		string ec_dp_dn_m_l_gain_pkt:source = "APID826:EC_DP_DN_M_L_GAIN_PKT" ;
  	ubyte ec_dp_hrd_pkt_norm_test(scans) ;
  		ec_dp_hrd_pkt_norm_test:_FillValue = 254UB ;
  		ec_dp_hrd_pkt_norm_test:valid_min = 0UB ;
  		ec_dp_hrd_pkt_norm_test:valid_max = 1UB ;
  		ec_dp_hrd_pkt_norm_test:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string ec_dp_hrd_pkt_norm_test:coordinates = "start_of_scan_time" ;
  		string ec_dp_hrd_pkt_norm_test:long_name = "Packet Normal/Test State" ;
  		string ec_dp_hrd_pkt_norm_test:source = "APID826:EC_DP_HRD_PKT_NORM_TEST" ;
  	ubyte ec_dp_nonrdt_fpie_pwr(scans) ;
  		ec_dp_nonrdt_fpie_pwr:_FillValue = 254UB ;
  		ec_dp_nonrdt_fpie_pwr:valid_min = 0UB ;
  		ec_dp_nonrdt_fpie_pwr:valid_max = 1UB ;
  		ec_dp_nonrdt_fpie_pwr:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string ec_dp_nonrdt_fpie_pwr:coordinates = "start_of_scan_time" ;
  		string ec_dp_nonrdt_fpie_pwr:long_name = "Non-redundant FPIE Power" ;
  		string ec_dp_nonrdt_fpie_pwr:source = "APID826:EC_DP_NONRDT_FPIE_PWR" ;
  	ubyte ec_dp_servo_in_use(scans) ;
  		ec_dp_servo_in_use:_FillValue = 254UB ;
  		ec_dp_servo_in_use:valid_min = 0UB ;
  		ec_dp_servo_in_use:valid_max = 1UB ;
  		ec_dp_servo_in_use:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string ec_dp_servo_in_use:coordinates = "start_of_scan_time" ;
  		string ec_dp_servo_in_use:long_name = "Servo In Use" ;
  		string ec_dp_servo_in_use:source = "APID826:EC_DP_SERVO_IN_USE" ;
  	ubyte ec_ps_sec_b_apfp_on(scans) ;
  		ec_ps_sec_b_apfp_on:_FillValue = 254UB ;
  		ec_ps_sec_b_apfp_on:valid_min = 0UB ;
  		ec_ps_sec_b_apfp_on:valid_max = 1UB ;
  		ec_ps_sec_b_apfp_on:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string ec_ps_sec_b_apfp_on:coordinates = "start_of_scan_time" ;
  		string ec_ps_sec_b_apfp_on:long_name = "Power Supply Section B ASP FPIE State" ;
  		string ec_ps_sec_b_apfp_on:source = "APID826:EC_PS_SEC_B_APFP_ON" ;
  	ubyte ec_ps_sec_c_se_on(scans) ;
  		ec_ps_sec_c_se_on:_FillValue = 254UB ;
  		ec_ps_sec_c_se_on:valid_min = 0UB ;
  		ec_ps_sec_c_se_on:valid_max = 1UB ;
  		ec_ps_sec_c_se_on:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string ec_ps_sec_c_se_on:coordinates = "start_of_scan_time" ;
  		string ec_ps_sec_c_se_on:long_name = "Power Supply Section C SCE State" ;
  		string ec_ps_sec_c_se_on:source = "APID826:EC_PS_SEC_C_SE_ON" ;
  	ubyte ec_ps_sec_d_csog_on(scans) ;
  		ec_ps_sec_d_csog_on:_FillValue = 254UB ;
  		ec_ps_sec_d_csog_on:valid_min = 0UB ;
  		ec_ps_sec_d_csog_on:valid_max = 1UB ;
  		ec_ps_sec_d_csog_on:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string ec_ps_sec_d_csog_on:coordinates = "start_of_scan_time" ;
  		string ec_ps_sec_d_csog_on:long_name = "Power Supply Section D Cold-Stage Outgas Heater State" ;
  		string ec_ps_sec_d_csog_on:source = "APID826:EC_PS_SEC_D_CSOG_ON" ;
  	ubyte ec_ps_sec_e_isog_on(scans) ;
  		ec_ps_sec_e_isog_on:_FillValue = 254UB ;
  		ec_ps_sec_e_isog_on:valid_min = 0UB ;
  		ec_ps_sec_e_isog_on:valid_max = 1UB ;
  		ec_ps_sec_e_isog_on:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string ec_ps_sec_e_isog_on:coordinates = "start_of_scan_time" ;
  		string ec_ps_sec_e_isog_on:long_name = "Power Supply Section E Intermediate-Stage Outgas Heater State" ;
  		string ec_ps_sec_e_isog_on:source = "APID826:EC_PS_SEC_E_ISOG_ON" ;
  	ubyte ec_se_a_anlg_pwr_on(scans) ;
  		ec_se_a_anlg_pwr_on:_FillValue = 254UB ;
  		ec_se_a_anlg_pwr_on:valid_min = 0UB ;
  		ec_se_a_anlg_pwr_on:valid_max = 1UB ;
  		ec_se_a_anlg_pwr_on:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string ec_se_a_anlg_pwr_on:coordinates = "start_of_scan_time" ;
  		string ec_se_a_anlg_pwr_on:long_name = "SCE-A Analog Power State" ;
  		string ec_se_a_anlg_pwr_on:source = "APID826:EC_SE_A_ANLG_PWR_ON" ;
  	ubyte ec_se_a_mtr_coil_driver(scans) ;
  		ec_se_a_mtr_coil_driver:_FillValue = 254UB ;
  		ec_se_a_mtr_coil_driver:valid_min = 0UB ;
  		ec_se_a_mtr_coil_driver:valid_max = 1UB ;
  		ec_se_a_mtr_coil_driver:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string ec_se_a_mtr_coil_driver:coordinates = "start_of_scan_time" ;
  		string ec_se_a_mtr_coil_driver:long_name = "SCE-A Motor Coil Driver Source" ;
  		string ec_se_a_mtr_coil_driver:source = "APID826:EC_SE_A_MTR_COIL_DRIVER" ;
  	ubyte ec_se_a_mtrs_stopped(scans) ;
  		ec_se_a_mtrs_stopped:_FillValue = 254UB ;
  		ec_se_a_mtrs_stopped:valid_min = 0UB ;
  		ec_se_a_mtrs_stopped:valid_max = 1UB ;
  		ec_se_a_mtrs_stopped:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string ec_se_a_mtrs_stopped:coordinates = "start_of_scan_time" ;
  		string ec_se_a_mtrs_stopped:long_name = "SCE-A Motor State" ;
  		string ec_se_a_mtrs_stopped:source = "APID826:EC_SE_A_MTRS_STOPPED" ;
  	ubyte ec_se_a_tele_pos_known(scans) ;
  		ec_se_a_tele_pos_known:_FillValue = 254UB ;
  		ec_se_a_tele_pos_known:valid_min = 0UB ;
  		ec_se_a_tele_pos_known:valid_max = 1UB ;
  		ec_se_a_tele_pos_known:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string ec_se_a_tele_pos_known:coordinates = "start_of_scan_time" ;
  		string ec_se_a_tele_pos_known:long_name = "SCE-A Telescope Position State" ;
  		string ec_se_a_tele_pos_known:source = "APID826:EC_SE_A_TELE_POS_KNOWN" ;
  	ubyte ec_se_b_anlg_pwr_on(scans) ;
  		ec_se_b_anlg_pwr_on:_FillValue = 254UB ;
  		ec_se_b_anlg_pwr_on:valid_min = 0UB ;
  		ec_se_b_anlg_pwr_on:valid_max = 1UB ;
  		ec_se_b_anlg_pwr_on:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string ec_se_b_anlg_pwr_on:coordinates = "start_of_scan_time" ;
  		string ec_se_b_anlg_pwr_on:long_name = "SCE-B Analog Power State" ;
  		string ec_se_b_anlg_pwr_on:source = "APID826:EC_SE_B_ANLG_PWR_ON" ;
  	ubyte ec_se_b_mtr_coil_driver(scans) ;
  		ec_se_b_mtr_coil_driver:_FillValue = 254UB ;
  		ec_se_b_mtr_coil_driver:valid_min = 0UB ;
  		ec_se_b_mtr_coil_driver:valid_max = 1UB ;
  		ec_se_b_mtr_coil_driver:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string ec_se_b_mtr_coil_driver:coordinates = "start_of_scan_time" ;
  		string ec_se_b_mtr_coil_driver:long_name = "SCE-B Motor Coil Driver Source" ;
  		string ec_se_b_mtr_coil_driver:source = "APID826:EC_SE_B_MTR_COIL_DRIVER" ;
  	ubyte ec_se_b_mtrs_stopped(scans) ;
  		ec_se_b_mtrs_stopped:_FillValue = 254UB ;
  		ec_se_b_mtrs_stopped:valid_min = 0UB ;
  		ec_se_b_mtrs_stopped:valid_max = 1UB ;
  		ec_se_b_mtrs_stopped:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string ec_se_b_mtrs_stopped:coordinates = "start_of_scan_time" ;
  		string ec_se_b_mtrs_stopped:long_name = "SCE-B Motor State" ;
  		string ec_se_b_mtrs_stopped:source = "APID826:EC_SE_B_MTRS_STOPPED" ;
  	ubyte ec_se_b_tele_pos_known(scans) ;
  		ec_se_b_tele_pos_known:_FillValue = 254UB ;
  		ec_se_b_tele_pos_known:valid_min = 0UB ;
  		ec_se_b_tele_pos_known:valid_max = 1UB ;
  		ec_se_b_tele_pos_known:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string ec_se_b_tele_pos_known:coordinates = "start_of_scan_time" ;
  		string ec_se_b_tele_pos_known:long_name = "SCE-B Telescope Position State" ;
  		string ec_se_b_tele_pos_known:source = "APID826:EC_SE_B_TELE_POS_KNOWN" ;
  	ubyte ec_dp_dn_aggreg_mode(scans) ;
  		ec_dp_dn_aggreg_mode:_FillValue = 254UB ;
  		ec_dp_dn_aggreg_mode:valid_min = 0UB ;
  		ec_dp_dn_aggreg_mode:valid_max = 63UB ;
  		ec_dp_dn_aggreg_mode:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string ec_dp_dn_aggreg_mode:coordinates = "start_of_scan_time" ;
  		string ec_dp_dn_aggreg_mode:long_name = "Day/Night Band Aggregation Mode" ;
  		string ec_dp_dn_aggreg_mode:source = "APID826:EC_DP_DN_AGGREG_MODE" ;
  	ubyte ec_cp_blk_pwr_sel(scans) ;
  		ec_cp_blk_pwr_sel:_FillValue = 254UB ;
  		ec_cp_blk_pwr_sel:valid_min = 0UB ;
  		ec_cp_blk_pwr_sel:valid_max = 1UB ;
  		ec_cp_blk_pwr_sel:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string ec_cp_blk_pwr_sel:coordinates = "start_of_scan_time" ;
  		string ec_cp_blk_pwr_sel:long_name = "Block Power Selection" ;
  		string ec_cp_blk_pwr_sel:source = "APID826:EC_CP_BLK_PWR_SEL" ;
  	ubyte ec_dp_ap_m16_tdi_on(scans) ;
  		ec_dp_ap_m16_tdi_on:_FillValue = 254UB ;
  		ec_dp_ap_m16_tdi_on:valid_min = 0UB ;
  		ec_dp_ap_m16_tdi_on:valid_max = 1UB ;
  		ec_dp_ap_m16_tdi_on:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string ec_dp_ap_m16_tdi_on:coordinates = "start_of_scan_time" ;
  		string ec_dp_ap_m16_tdi_on:long_name = "ASP M16 Time Delay Integration State" ;
  		string ec_dp_ap_m16_tdi_on:source = "APID826:EC_DP_AP_M16_TDI_ON" ;
  	ushort ec_dp_scan_encdr_delta(scans) ;
  		ec_dp_scan_encdr_delta:_FillValue = 65534US ;
  		ec_dp_scan_encdr_delta:valid_min = 0US ;
  		ec_dp_scan_encdr_delta:valid_max = 32767US ;
  		ec_dp_scan_encdr_delta:missing_value = 65528US, 65529US, 65530US, 65531US, 65532US, 65533US, 65534US, 65535US ;
  		string ec_dp_scan_encdr_delta:coordinates = "start_of_scan_time" ;
  		string ec_dp_scan_encdr_delta:long_name = "Scan Encoder Delta" ;
  		string ec_dp_scan_encdr_delta:source = "APID826:EC_DP_SCAN_ENCDR_DELTA" ;
  	ubyte ec_dp_ap_self_test(scans) ;
  		ec_dp_ap_self_test:_FillValue = 254UB ;
  		ec_dp_ap_self_test:valid_min = 0UB ;
  		ec_dp_ap_self_test:valid_max = 1UB ;
  		ec_dp_ap_self_test:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string ec_dp_ap_self_test:coordinates = "start_of_scan_time" ;
  		string ec_dp_ap_self_test:long_name = "Self-test State" ;
  		string ec_dp_ap_self_test:source = "APID826:EC_DP_AP_SELF_TEST" ;
  	ubyte ec_se_servo_pwr_sel(scans) ;
  		ec_se_servo_pwr_sel:_FillValue = 254UB ;
  		ec_se_servo_pwr_sel:valid_min = 0UB ;
  		ec_se_servo_pwr_sel:valid_max = 1UB ;
  		ec_se_servo_pwr_sel:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string ec_se_servo_pwr_sel:coordinates = "start_of_scan_time" ;
  		string ec_se_servo_pwr_sel:long_name = "SCE Servo Power Selection" ;
  		string ec_se_servo_pwr_sel:source = "APID826:EC_SE_SERVO_PWR_SEL" ;
  	ubyte ec_dp_dnb_1a_1b_stage(scans) ;
  		ec_dp_dnb_1a_1b_stage:_FillValue = 254UB ;
  		ec_dp_dnb_1a_1b_stage:valid_min = 0UB ;
  		ec_dp_dnb_1a_1b_stage:valid_max = 2UB ;
  		ec_dp_dnb_1a_1b_stage:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string ec_dp_dnb_1a_1b_stage:coordinates = "start_of_scan_time" ;
  		string ec_dp_dnb_1a_1b_stage:long_name = "Day/Night Band Stage 1 Data Selection" ;
  		string ec_dp_dnb_1a_1b_stage:source = "APID826:EC_DP_DNB_1A_1B_STAGE" ;
  	ubyte ec_dp_dnb_tmg_mode(scans) ;
  		ec_dp_dnb_tmg_mode:_FillValue = 254UB ;
  		ec_dp_dnb_tmg_mode:valid_min = 0UB ;
  		ec_dp_dnb_tmg_mode:valid_max = 1UB ;
  		ec_dp_dnb_tmg_mode:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string ec_dp_dnb_tmg_mode:coordinates = "start_of_scan_time" ;
  		string ec_dp_dnb_tmg_mode:long_name = "Day/Night Band Timing Mode" ;
  		string ec_dp_dnb_tmg_mode:source = "APID826:EC_DP_DNB_TMG_MODE" ;
  	ubyte ec_dp_dnb_dark_sub_cal(scans) ;
  		ec_dp_dnb_dark_sub_cal:_FillValue = 254UB ;
  		ec_dp_dnb_dark_sub_cal:valid_min = 0UB ;
  		ec_dp_dnb_dark_sub_cal:valid_max = 1UB ;
  		ec_dp_dnb_dark_sub_cal:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string ec_dp_dnb_dark_sub_cal:coordinates = "start_of_scan_time" ;
  		string ec_dp_dnb_dark_sub_cal:long_name = "Day/Night Band Calibview Dark Pixel Subtraction" ;
  		string ec_dp_dnb_dark_sub_cal:source = "APID826:EC_DP_DNB_DARK_SUB_CAL" ;
  	ubyte ec_dp_dnb_dark_sub_eth(scans) ;
  		ec_dp_dnb_dark_sub_eth:_FillValue = 254UB ;
  		ec_dp_dnb_dark_sub_eth:valid_min = 0UB ;
  		ec_dp_dnb_dark_sub_eth:valid_max = 1UB ;
  		ec_dp_dnb_dark_sub_eth:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string ec_dp_dnb_dark_sub_eth:coordinates = "start_of_scan_time" ;
  		string ec_dp_dnb_dark_sub_eth:long_name = "Day/Night Band Earthview Dark Pixel Subtraction" ;
  		string ec_dp_dnb_dark_sub_eth:source = "APID826:EC_DP_DNB_DARK_SUB_ETH" ;
  	ubyte ec_ap_dc_fast_restore(scans) ;
  		ec_ap_dc_fast_restore:_FillValue = 254UB ;
  		ec_ap_dc_fast_restore:valid_min = 0UB ;
  		ec_ap_dc_fast_restore:valid_max = 1UB ;
  		ec_ap_dc_fast_restore:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string ec_ap_dc_fast_restore:coordinates = "start_of_scan_time" ;
  		string ec_ap_dc_fast_restore:long_name = "ASP Restore Algorithm" ;
  		string ec_ap_dc_fast_restore:source = "APID826:EC_AP_DC_FAST_RESTORE" ;
  	ubyte es_se_a_ham_mir_side(scans) ;
  		es_se_a_ham_mir_side:_FillValue = 254UB ;
  		es_se_a_ham_mir_side:valid_min = 0UB ;
  		es_se_a_ham_mir_side:valid_max = 1UB ;
  		es_se_a_ham_mir_side:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string es_se_a_ham_mir_side:coordinates = "start_of_scan_time" ;
  		string es_se_a_ham_mir_side:long_name = "SCE-A Half-Angle Mirror Side" ;
  		string es_se_a_ham_mir_side:source = "APID826:ES_SE_A_HAM_MIR_SIDE" ;
  	ubyte es_se_b_ham_mir_side(scans) ;
  		es_se_b_ham_mir_side:_FillValue = 254UB ;
  		es_se_b_ham_mir_side:valid_min = 0UB ;
  		es_se_b_ham_mir_side:valid_max = 1UB ;
  		es_se_b_ham_mir_side:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string es_se_b_ham_mir_side:coordinates = "start_of_scan_time" ;
  		string es_se_b_ham_mir_side:long_name = "SCE-B Half-Angle Mirror Side" ;
  		string es_se_b_ham_mir_side:source = "APID826:ES_SE_B_HAM_MIR_SIDE" ;
  	short ei_se_a_ham_mtr_curr(scans) ;
  		ei_se_a_ham_mtr_curr:_FillValue = -998s ;
  		ei_se_a_ham_mtr_curr:valid_min = -8192s ;
  		ei_se_a_ham_mtr_curr:valid_max = 8191s ;
  		ei_se_a_ham_mtr_curr:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string ei_se_a_ham_mtr_curr:coordinates = "start_of_scan_time" ;
  		string ei_se_a_ham_mtr_curr:long_name = "SCE-A Half-Angle Mirror Motor Current" ;
  		string ei_se_a_ham_mtr_curr:source = "APID826:EI_SE_A_HAM_MTR_CURR" ;
  	short ei_se_a_tele_mtr_curr(scans) ;
  		ei_se_a_tele_mtr_curr:_FillValue = -998s ;
  		ei_se_a_tele_mtr_curr:valid_min = -8192s ;
  		ei_se_a_tele_mtr_curr:valid_max = 8191s ;
  		ei_se_a_tele_mtr_curr:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string ei_se_a_tele_mtr_curr:coordinates = "start_of_scan_time" ;
  		string ei_se_a_tele_mtr_curr:long_name = "SCE-A Telescope Motor Current" ;
  		string ei_se_a_tele_mtr_curr:source = "APID826:EI_SE_A_TELE_MTR_CURR" ;
  	short ei_se_b_ham_mtr_curr(scans) ;
  		ei_se_b_ham_mtr_curr:_FillValue = -998s ;
  		ei_se_b_ham_mtr_curr:valid_min = -8192s ;
  		ei_se_b_ham_mtr_curr:valid_max = 8191s ;
  		ei_se_b_ham_mtr_curr:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string ei_se_b_ham_mtr_curr:coordinates = "start_of_scan_time" ;
  		string ei_se_b_ham_mtr_curr:long_name = "SCE-B Half-Angle Mirror Motor Current" ;
  		string ei_se_b_ham_mtr_curr:source = "APID826:EI_SE_B_HAM_MTR_CURR" ;
  	short ei_se_b_tele_mtr_curr(scans) ;
  		ei_se_b_tele_mtr_curr:_FillValue = -998s ;
  		ei_se_b_tele_mtr_curr:valid_min = -8192s ;
  		ei_se_b_tele_mtr_curr:valid_max = 8191s ;
  		ei_se_b_tele_mtr_curr:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string ei_se_b_tele_mtr_curr:coordinates = "start_of_scan_time" ;
  		string ei_se_b_tele_mtr_curr:long_name = "SCE-B Telescope Motor Current" ;
  		string ei_se_b_tele_mtr_curr:source = "APID826:EI_SE_B_TELE_MTR_CURR" ;
  	short ev_ct_prec_tref_mux1ca1(scans) ;
  		ev_ct_prec_tref_mux1ca1:_FillValue = -998s ;
  		ev_ct_prec_tref_mux1ca1:valid_min = -8192s ;
  		ev_ct_prec_tref_mux1ca1:valid_max = 8191s ;
  		ev_ct_prec_tref_mux1ca1:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string ev_ct_prec_tref_mux1ca1:coordinates = "start_of_scan_time" ;
  		string ev_ct_prec_tref_mux1ca1:long_name = "Precision Calibration Reference Thermistor Mux1Cal1 Voltage" ;
  		string ev_ct_prec_tref_mux1ca1:source = "APID826:EV_CT_PREC_TREF_MUX1CA1" ;
  	short ev_ct_prec_tref_mux1ca2(scans) ;
  		ev_ct_prec_tref_mux1ca2:_FillValue = -998s ;
  		ev_ct_prec_tref_mux1ca2:valid_min = -8192s ;
  		ev_ct_prec_tref_mux1ca2:valid_max = 8191s ;
  		ev_ct_prec_tref_mux1ca2:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string ev_ct_prec_tref_mux1ca2:coordinates = "start_of_scan_time" ;
  		string ev_ct_prec_tref_mux1ca2:long_name = "Precision Calibration Reference Thermistor Mux1Cal2 Voltage" ;
  		string ev_ct_prec_tref_mux1ca2:source = "APID826:EV_CT_PREC_TREF_MUX1CA2" ;
  	short ev_ct_prec_tref_mux1ca3(scans) ;
  		ev_ct_prec_tref_mux1ca3:_FillValue = -998s ;
  		ev_ct_prec_tref_mux1ca3:valid_min = -8192s ;
  		ev_ct_prec_tref_mux1ca3:valid_max = 8191s ;
  		ev_ct_prec_tref_mux1ca3:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string ev_ct_prec_tref_mux1ca3:coordinates = "start_of_scan_time" ;
  		string ev_ct_prec_tref_mux1ca3:long_name = "Precision Calibration Reference Thermistor Mux1Cal3 Voltage" ;
  		string ev_ct_prec_tref_mux1ca3:source = "APID826:EV_CT_PREC_TREF_MUX1CA3" ;
  	short ev_ft_adc_ref(scans) ;
  		ev_ft_adc_ref:_FillValue = -998s ;
  		ev_ft_adc_ref:valid_min = -8192s ;
  		ev_ft_adc_ref:valid_max = 8191s ;
  		ev_ft_adc_ref:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string ev_ft_adc_ref:coordinates = "start_of_scan_time" ;
  		string ev_ft_adc_ref:long_name = "FTC ADC 5 Volt Reference Voltage" ;
  		string ev_ft_adc_ref:source = "APID826:EV_FT_ADC_REF" ;
  	short ev_ft_adc_ref_lw_stpt(scans) ;
  		ev_ft_adc_ref_lw_stpt:_FillValue = -998s ;
  		ev_ft_adc_ref_lw_stpt:valid_min = -8192s ;
  		ev_ft_adc_ref_lw_stpt:valid_max = 8191s ;
  		ev_ft_adc_ref_lw_stpt:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string ev_ft_adc_ref_lw_stpt:coordinates = "start_of_scan_time" ;
  		string ev_ft_adc_ref_lw_stpt:long_name = "FTC ADC Long-Wavelength Setpoint Reference Voltage" ;
  		string ev_ft_adc_ref_lw_stpt:source = "APID826:EV_FT_ADC_REF_LW_STPT" ;
  	short ev_ft_ckt_gnd(scans) ;
  		ev_ft_ckt_gnd:_FillValue = -998s ;
  		ev_ft_ckt_gnd:valid_min = -8192s ;
  		ev_ft_ckt_gnd:valid_max = 8191s ;
  		ev_ft_ckt_gnd:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string ev_ft_ckt_gnd:coordinates = "start_of_scan_time" ;
  		string ev_ft_ckt_gnd:long_name = "FTC Circuit Ground Voltage" ;
  		string ev_ft_ckt_gnd:source = "APID826:EV_FT_CKT_GND" ;
  	short ev_ft_lw_cfpa_htr_pwr(scans) ;
  		ev_ft_lw_cfpa_htr_pwr:_FillValue = -998s ;
  		ev_ft_lw_cfpa_htr_pwr:valid_min = -8192s ;
  		ev_ft_lw_cfpa_htr_pwr:valid_max = 8191s ;
  		ev_ft_lw_cfpa_htr_pwr:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string ev_ft_lw_cfpa_htr_pwr:coordinates = "start_of_scan_time" ;
  		string ev_ft_lw_cfpa_htr_pwr:long_name = "FTC Long-WavelengthFPA Heater Power Supply Voltage" ;
  		string ev_ft_lw_cfpa_htr_pwr:source = "APID826:EV_FT_LW_CFPA_HTR_PWR" ;
  	short ev_ft_lw_setpt_ref(scans) ;
  		ev_ft_lw_setpt_ref:_FillValue = -998s ;
  		ev_ft_lw_setpt_ref:valid_min = -8192s ;
  		ev_ft_lw_setpt_ref:valid_max = 8191s ;
  		ev_ft_lw_setpt_ref:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string ev_ft_lw_setpt_ref:coordinates = "start_of_scan_time" ;
  		string ev_ft_lw_setpt_ref:long_name = "FTC Long-Wavelength Setpoint Reference Voltage" ;
  		string ev_ft_lw_setpt_ref:source = "APID826:EV_FT_LW_SETPT_REF" ;
  	short ev_ft_sm_cfpa_htr_pwr(scans) ;
  		ev_ft_sm_cfpa_htr_pwr:_FillValue = -998s ;
  		ev_ft_sm_cfpa_htr_pwr:valid_min = -8192s ;
  		ev_ft_sm_cfpa_htr_pwr:valid_max = 8191s ;
  		ev_ft_sm_cfpa_htr_pwr:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string ev_ft_sm_cfpa_htr_pwr:coordinates = "start_of_scan_time" ;
  		string ev_ft_sm_cfpa_htr_pwr:long_name = "FTC Short/Medium-Wavelength FPA Heater Power Supply Voltage" ;
  		string ev_ft_sm_cfpa_htr_pwr:source = "APID826:EV_FT_SM_CFPA_HTR_PWR" ;
  	short ev_ft_sm_setpt_ref(scans) ;
  		ev_ft_sm_setpt_ref:_FillValue = -998s ;
  		ev_ft_sm_setpt_ref:valid_min = -8192s ;
  		ev_ft_sm_setpt_ref:valid_max = 8191s ;
  		ev_ft_sm_setpt_ref:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string ev_ft_sm_setpt_ref:coordinates = "start_of_scan_time" ;
  		string ev_ft_sm_setpt_ref:long_name = "FTC Short/Medium-Wavelength Setpoint Reference Voltage" ;
  		string ev_ft_sm_setpt_ref:source = "APID826:EV_FT_SM_SETPT_REF" ;
  	short ev_se_a_ham_rate_error(scans) ;
  		ev_se_a_ham_rate_error:_FillValue = -998s ;
  		ev_se_a_ham_rate_error:valid_min = -8192s ;
  		ev_se_a_ham_rate_error:valid_max = 8191s ;
  		ev_se_a_ham_rate_error:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string ev_se_a_ham_rate_error:coordinates = "start_of_scan_time" ;
  		string ev_se_a_ham_rate_error:long_name = "SCE-A Half-Angle Mirror Rate Error Voltage" ;
  		string ev_se_a_ham_rate_error:source = "APID826:EV_SE_A_HAM_RATE_ERROR" ;
  	short ev_se_a_tele_rate_error(scans) ;
  		ev_se_a_tele_rate_error:_FillValue = -998s ;
  		ev_se_a_tele_rate_error:valid_min = -8192s ;
  		ev_se_a_tele_rate_error:valid_max = 8191s ;
  		ev_se_a_tele_rate_error:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string ev_se_a_tele_rate_error:coordinates = "start_of_scan_time" ;
  		string ev_se_a_tele_rate_error:long_name = "SCE-A Telescope Rate Error Voltage" ;
  		string ev_se_a_tele_rate_error:source = "APID826:EV_SE_A_TELE_RATE_ERROR" ;
  	short ev_se_b_ham_rate_error(scans) ;
  		ev_se_b_ham_rate_error:_FillValue = -998s ;
  		ev_se_b_ham_rate_error:valid_min = -8192s ;
  		ev_se_b_ham_rate_error:valid_max = 8191s ;
  		ev_se_b_ham_rate_error:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string ev_se_b_ham_rate_error:coordinates = "start_of_scan_time" ;
  		string ev_se_b_ham_rate_error:long_name = "SCE-B Half-Angle Mirror Rate Error Voltage" ;
  		string ev_se_b_ham_rate_error:source = "APID826:EV_SE_B_HAM_RATE_ERROR" ;
  	short ev_se_b_tele_rate_error(scans) ;
  		ev_se_b_tele_rate_error:_FillValue = -998s ;
  		ev_se_b_tele_rate_error:valid_min = -8192s ;
  		ev_se_b_tele_rate_error:valid_max = 8191s ;
  		ev_se_b_tele_rate_error:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string ev_se_b_tele_rate_error:coordinates = "start_of_scan_time" ;
  		string ev_se_b_tele_rate_error:long_name = "SCE-B Telescope Rate Error Voltage" ;
  		string ev_se_b_tele_rate_error:source = "APID826:EV_SE_B_TELE_RATE_ERROR" ;
  	ubyte c_ap_visnir_reg_tbl_rev(scans) ;
  		c_ap_visnir_reg_tbl_rev:_FillValue = 254UB ;
  		c_ap_visnir_reg_tbl_rev:valid_min = 0UB ;
  		c_ap_visnir_reg_tbl_rev:valid_max = 248UB ;
  		c_ap_visnir_reg_tbl_rev:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string c_ap_visnir_reg_tbl_rev:coordinates = "start_of_scan_time" ;
  		string c_ap_visnir_reg_tbl_rev:long_name = "ASP Visible/NIR Register Table Revision" ;
  		string c_ap_visnir_reg_tbl_rev:source = "APID826:C_AP_VISNIR_REG_TBL_REV" ;
  	ubyte c_ap_smwir_reg_tbl_rev(scans) ;
  		c_ap_smwir_reg_tbl_rev:_FillValue = 254UB ;
  		c_ap_smwir_reg_tbl_rev:valid_min = 0UB ;
  		c_ap_smwir_reg_tbl_rev:valid_max = 248UB ;
  		c_ap_smwir_reg_tbl_rev:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string c_ap_smwir_reg_tbl_rev:coordinates = "start_of_scan_time" ;
  		string c_ap_smwir_reg_tbl_rev:long_name = "ASP SW/MW-IR Register Table Revision" ;
  		string c_ap_smwir_reg_tbl_rev:source = "APID826:C_AP_SMWIR_REG_TBL_REV" ;
  	ubyte c_ap_lwir_reg_tbl_rev(scans) ;
  		c_ap_lwir_reg_tbl_rev:_FillValue = 254UB ;
  		c_ap_lwir_reg_tbl_rev:valid_min = 0UB ;
  		c_ap_lwir_reg_tbl_rev:valid_max = 248UB ;
  		c_ap_lwir_reg_tbl_rev:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string c_ap_lwir_reg_tbl_rev:coordinates = "start_of_scan_time" ;
  		string c_ap_lwir_reg_tbl_rev:long_name = "ASP LW-IR Register Table Revision" ;
  		string c_ap_lwir_reg_tbl_rev:source = "APID826:C_AP_LWIR_REG_TBL_REV" ;
  	ubyte c_ap_fpa_ideal_tbl_rev(scans) ;
  		c_ap_fpa_ideal_tbl_rev:_FillValue = 254UB ;
  		c_ap_fpa_ideal_tbl_rev:valid_min = 0UB ;
  		c_ap_fpa_ideal_tbl_rev:valid_max = 248UB ;
  		c_ap_fpa_ideal_tbl_rev:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string c_ap_fpa_ideal_tbl_rev:coordinates = "start_of_scan_time" ;
  		string c_ap_fpa_ideal_tbl_rev:long_name = "ASP FPA Ideal Offsets Table Revision" ;
  		string c_ap_fpa_ideal_tbl_rev:source = "APID826:C_AP_FPA_IDEAL_TBL_REV" ;
  	ubyte ec_ap_dc_restore(scans) ;
  		ec_ap_dc_restore:_FillValue = 254UB ;
  		ec_ap_dc_restore:valid_min = 0UB ;
  		ec_ap_dc_restore:valid_max = 1UB ;
  		ec_ap_dc_restore:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string ec_ap_dc_restore:coordinates = "start_of_scan_time" ;
  		string ec_ap_dc_restore:long_name = "ASP Global DC Restore State" ;
  		string ec_ap_dc_restore:source = "APID826:EC_AP_DC_RESTORE" ;
  	ubyte ec_ap_det_connected(scans) ;
  		ec_ap_det_connected:_FillValue = 254UB ;
  		ec_ap_det_connected:valid_min = 0UB ;
  		ec_ap_det_connected:valid_max = 1UB ;
  		ec_ap_det_connected:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string ec_ap_det_connected:coordinates = "start_of_scan_time" ;
  		string ec_ap_det_connected:long_name = "ASP Detector State" ;
  		string ec_ap_det_connected:source = "APID826:EC_AP_DET_CONNECTED" ;
  	ubyte ec_ap_lw_ifs_width(scans) ;
  		ec_ap_lw_ifs_width:_FillValue = 254UB ;
  		ec_ap_lw_ifs_width:valid_min = 2UB ;
  		ec_ap_lw_ifs_width:valid_max = 16UB ;
  		ec_ap_lw_ifs_width:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string ec_ap_lw_ifs_width:coordinates = "start_of_scan_time" ;
  		string ec_ap_lw_ifs_width:units = "ticks" ;
  		string ec_ap_lw_ifs_width:long_name = "ASP LW-IR Imaging Frame Sync Width" ;
  		string ec_ap_lw_ifs_width:source = "APID826:EC_AP_LW_IFS_WIDTH" ;
  	ubyte ec_ap_dual_gain_3_ops(scans) ;
  		ec_ap_dual_gain_3_ops:_FillValue = 254UB ;
  		ec_ap_dual_gain_3_ops:valid_min = 0UB ;
  		ec_ap_dual_gain_3_ops:valid_max = 2UB ;
  		ec_ap_dual_gain_3_ops:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string ec_ap_dual_gain_3_ops:coordinates = "start_of_scan_time" ;
  		string ec_ap_dual_gain_3_ops:long_name = "ASP Dual Gain Operation Mode" ;
  		string ec_ap_dual_gain_3_ops:source = "APID826:EC_AP_DUAL_GAIN_3_OPS" ;
  	ubyte ec_ap_lw_rfs_width(scans) ;
  		ec_ap_lw_rfs_width:_FillValue = 254UB ;
  		ec_ap_lw_rfs_width:valid_min = 2UB ;
  		ec_ap_lw_rfs_width:valid_max = 36UB ;
  		ec_ap_lw_rfs_width:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string ec_ap_lw_rfs_width:coordinates = "start_of_scan_time" ;
  		string ec_ap_lw_rfs_width:units = "ticks" ;
  		string ec_ap_lw_rfs_width:long_name = "ASP LW-IR Radiometric Frame Sync Width" ;
  		string ec_ap_lw_rfs_width:source = "APID826:EC_AP_LW_RFS_WIDTH" ;
  	ubyte ec_ap_fpa_st_3_ops(scans) ;
  		ec_ap_fpa_st_3_ops:_FillValue = 254UB ;
  		ec_ap_fpa_st_3_ops:valid_min = 0UB ;
  		ec_ap_fpa_st_3_ops:valid_max = 2UB ;
  		ec_ap_fpa_st_3_ops:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string ec_ap_fpa_st_3_ops:coordinates = "start_of_scan_time" ;
  		string ec_ap_fpa_st_3_ops:long_name = "ASP FPA Self-test Operation Mode" ;
  		string ec_ap_fpa_st_3_ops:source = "APID826:EC_AP_FPA_ST_3_OPS" ;
  	ubyte ec_ap_sm_ifs_width(scans) ;
  		ec_ap_sm_ifs_width:_FillValue = 254UB ;
  		ec_ap_sm_ifs_width:valid_min = 2UB ;
  		ec_ap_sm_ifs_width:valid_max = 15UB ;
  		ec_ap_sm_ifs_width:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string ec_ap_sm_ifs_width:coordinates = "start_of_scan_time" ;
  		string ec_ap_sm_ifs_width:units = "ticks" ;
  		string ec_ap_sm_ifs_width:long_name = "ASP SW/MW-IR Imaging Frame Sync Width" ;
  		string ec_ap_sm_ifs_width:source = "APID826:EC_AP_SM_IFS_WIDTH" ;
  	ubyte ec_ap_sm_rfs_width(scans) ;
  		ec_ap_sm_rfs_width:_FillValue = 254UB ;
  		ec_ap_sm_rfs_width:valid_min = 2UB ;
  		ec_ap_sm_rfs_width:valid_max = 35UB ;
  		ec_ap_sm_rfs_width:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string ec_ap_sm_rfs_width:coordinates = "start_of_scan_time" ;
  		string ec_ap_sm_rfs_width:units = "ticks" ;
  		string ec_ap_sm_rfs_width:long_name = "ASP SW/MW-IR Radiometric Frame Sync Width" ;
  		string ec_ap_sm_rfs_width:source = "APID826:EC_AP_SM_RFS_WIDTH" ;
  	ubyte ec_ap_vn_ifs_width(scans) ;
  		ec_ap_vn_ifs_width:_FillValue = 254UB ;
  		ec_ap_vn_ifs_width:valid_min = 2UB ;
  		ec_ap_vn_ifs_width:valid_max = 15UB ;
  		ec_ap_vn_ifs_width:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string ec_ap_vn_ifs_width:coordinates = "start_of_scan_time" ;
  		string ec_ap_vn_ifs_width:units = "ticks" ;
  		string ec_ap_vn_ifs_width:long_name = "ASP Visible/NIR Imaging Frame Sync Width" ;
  		string ec_ap_vn_ifs_width:source = "APID826:EC_AP_VN_IFS_WIDTH" ;
  	ubyte ec_ap_vn_rfs_width(scans) ;
  		ec_ap_vn_rfs_width:_FillValue = 254UB ;
  		ec_ap_vn_rfs_width:valid_min = 2UB ;
  		ec_ap_vn_rfs_width:valid_max = 35UB ;
  		ec_ap_vn_rfs_width:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string ec_ap_vn_rfs_width:coordinates = "start_of_scan_time" ;
  		string ec_ap_vn_rfs_width:units = "ticks" ;
  		string ec_ap_vn_rfs_width:long_name = "ASP Visible/NIR Radiometric Frame Sync Width" ;
  		string ec_ap_vn_rfs_width:source = "APID826:EC_AP_VN_RFS_WIDTH" ;
  	short eta_ft_lw_cfpa_hi_rsl(scans) ;
  		eta_ft_lw_cfpa_hi_rsl:_FillValue = -998s ;
  		eta_ft_lw_cfpa_hi_rsl:valid_min = -8192s ;
  		eta_ft_lw_cfpa_hi_rsl:valid_max = 8191s ;
  		eta_ft_lw_cfpa_hi_rsl:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string eta_ft_lw_cfpa_hi_rsl:coordinates = "start_of_scan_time" ;
  		string eta_ft_lw_cfpa_hi_rsl:long_name = "LW-IR Cold FPA High Resolution Temperature" ;
  		string eta_ft_lw_cfpa_hi_rsl:source = "APID826:ETA_FT_LW_CFPA_HI_RSL" ;
  	short eta_ft_lw_cfpa_lo_rsl(scans) ;
  		eta_ft_lw_cfpa_lo_rsl:_FillValue = -998s ;
  		eta_ft_lw_cfpa_lo_rsl:valid_min = -8192s ;
  		eta_ft_lw_cfpa_lo_rsl:valid_max = 8191s ;
  		eta_ft_lw_cfpa_lo_rsl:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string eta_ft_lw_cfpa_lo_rsl:coordinates = "start_of_scan_time" ;
  		string eta_ft_lw_cfpa_lo_rsl:long_name = "LW-IR Cold FPA Low Resolution Temperature" ;
  		string eta_ft_lw_cfpa_lo_rsl:source = "APID826:ETA_FT_LW_CFPA_LO_RSL" ;
  	short eta_ft_sm_cfpa_hi_rsl(scans) ;
  		eta_ft_sm_cfpa_hi_rsl:_FillValue = -998s ;
  		eta_ft_sm_cfpa_hi_rsl:valid_min = -8192s ;
  		eta_ft_sm_cfpa_hi_rsl:valid_max = 8191s ;
  		eta_ft_sm_cfpa_hi_rsl:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string eta_ft_sm_cfpa_hi_rsl:coordinates = "start_of_scan_time" ;
  		string eta_ft_sm_cfpa_hi_rsl:long_name = "SW/MW-IR Cold FPA High Resolution Temperature" ;
  		string eta_ft_sm_cfpa_hi_rsl:source = "APID826:ETA_FT_SM_CFPA_HI_RSL" ;
  	short eta_ft_sm_cfpa_lo_rsl(scans) ;
  		eta_ft_sm_cfpa_lo_rsl:_FillValue = -998s ;
  		eta_ft_sm_cfpa_lo_rsl:valid_min = -8192s ;
  		eta_ft_sm_cfpa_lo_rsl:valid_max = 8191s ;
  		eta_ft_sm_cfpa_lo_rsl:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string eta_ft_sm_cfpa_lo_rsl:coordinates = "start_of_scan_time" ;
  		string eta_ft_sm_cfpa_lo_rsl:long_name = "SW/MW-IR Cold FPA Low Resolution Temperature" ;
  		string eta_ft_sm_cfpa_lo_rsl:source = "APID826:ETA_FT_SM_CFPA_LO_RSL" ;
  	short eta_ft_vis_nir_fpa(scans) ;
  		eta_ft_vis_nir_fpa:_FillValue = -998s ;
  		eta_ft_vis_nir_fpa:valid_min = -8192s ;
  		eta_ft_vis_nir_fpa:valid_max = 8191s ;
  		eta_ft_vis_nir_fpa:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string eta_ft_vis_nir_fpa:coordinates = "start_of_scan_time" ;
  		string eta_ft_vis_nir_fpa:long_name = "Visible/NIR FPA Temperature" ;
  		string eta_ft_vis_nir_fpa:source = "APID826:ETA_FT_VIS_NIR_FPA" ;
  	ubyte c_dp_aggreg_mode_rev(scans) ;
  		c_dp_aggreg_mode_rev:_FillValue = 254UB ;
  		c_dp_aggreg_mode_rev:valid_min = 0UB ;
  		c_dp_aggreg_mode_rev:valid_max = 248UB ;
  		c_dp_aggreg_mode_rev:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string c_dp_aggreg_mode_rev:coordinates = "start_of_scan_time" ;
  		string c_dp_aggreg_mode_rev:long_name = "Day/Night Band Aggregation Mode Revision" ;
  		string c_dp_aggreg_mode_rev:source = "APID826:C_DP_AGGREG_MODE_REV" ;
  	ubyte c_dp_threshold_tbl_rev(scans) ;
  		c_dp_threshold_tbl_rev:_FillValue = 254UB ;
  		c_dp_threshold_tbl_rev:valid_min = 0UB ;
  		c_dp_threshold_tbl_rev:valid_max = 248UB ;
  		c_dp_threshold_tbl_rev:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string c_dp_threshold_tbl_rev:coordinates = "start_of_scan_time" ;
  		string c_dp_threshold_tbl_rev:long_name = "Day/Night Band Threshold Table Revision" ;
  		string c_dp_threshold_tbl_rev:source = "APID826:C_DP_THRESHOLD_TBL_REV" ;
  	ubyte c_dp_1a_offsets_tbl_rev(scans) ;
  		c_dp_1a_offsets_tbl_rev:_FillValue = 254UB ;
  		c_dp_1a_offsets_tbl_rev:valid_min = 0UB ;
  		c_dp_1a_offsets_tbl_rev:valid_max = 248UB ;
  		c_dp_1a_offsets_tbl_rev:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string c_dp_1a_offsets_tbl_rev:coordinates = "start_of_scan_time" ;
  		string c_dp_1a_offsets_tbl_rev:long_name = "Day/Night Band 1A Offsets Table Revision" ;
  		string c_dp_1a_offsets_tbl_rev:source = "APID826:C_DP_1A_OFFSETS_TBL_REV" ;
  	short eta_dp_dnb_ccd(scans) ;
  		eta_dp_dnb_ccd:_FillValue = -998s ;
  		eta_dp_dnb_ccd:valid_min = -8192s ;
  		eta_dp_dnb_ccd:valid_max = 8191s ;
  		eta_dp_dnb_ccd:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string eta_dp_dnb_ccd:coordinates = "start_of_scan_time" ;
  		string eta_dp_dnb_ccd:long_name = "Day/Night Band CCD Temperature" ;
  		string eta_dp_dnb_ccd:source = "APID826:ETA_DP_DNB_CCD" ;
  	ubyte c_dp_1b_offsets_tbl_rev(scans) ;
  		c_dp_1b_offsets_tbl_rev:_FillValue = 254UB ;
  		c_dp_1b_offsets_tbl_rev:valid_min = 0UB ;
  		c_dp_1b_offsets_tbl_rev:valid_max = 248UB ;
  		c_dp_1b_offsets_tbl_rev:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string c_dp_1b_offsets_tbl_rev:coordinates = "start_of_scan_time" ;
  		string c_dp_1b_offsets_tbl_rev:long_name = "Day/Night Band 1B Offsets Table Revision" ;
  		string c_dp_1b_offsets_tbl_rev:source = "APID826:C_DP_1B_OFFSETS_TBL_REV" ;
  	ubyte c_dp_2_offsets_tbl_rev(scans) ;
  		c_dp_2_offsets_tbl_rev:_FillValue = 254UB ;
  		c_dp_2_offsets_tbl_rev:valid_min = 0UB ;
  		c_dp_2_offsets_tbl_rev:valid_max = 248UB ;
  		c_dp_2_offsets_tbl_rev:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string c_dp_2_offsets_tbl_rev:coordinates = "start_of_scan_time" ;
  		string c_dp_2_offsets_tbl_rev:long_name = "Day/Night Band 2 Offsets Table Revision" ;
  		string c_dp_2_offsets_tbl_rev:source = "APID826:C_DP_2_OFFSETS_TBL_REV" ;
  	ubyte c_dp_3_offsets_tbl_rev(scans) ;
  		c_dp_3_offsets_tbl_rev:_FillValue = 254UB ;
  		c_dp_3_offsets_tbl_rev:valid_min = 0UB ;
  		c_dp_3_offsets_tbl_rev:valid_max = 248UB ;
  		c_dp_3_offsets_tbl_rev:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string c_dp_3_offsets_tbl_rev:coordinates = "start_of_scan_time" ;
  		string c_dp_3_offsets_tbl_rev:long_name = "Day/Night Band 3 Offsets Table Revision" ;
  		string c_dp_3_offsets_tbl_rev:source = "APID826:C_DP_3_OFFSETS_TBL_REV" ;
  	ushort c_ap_m1_offsets(scans, mirror_sides, detectors_750m) ;
  		c_ap_m1_offsets:_FillValue = 65534US ;
  		c_ap_m1_offsets:valid_min = 0US ;
  		c_ap_m1_offsets:valid_max = 65535US ;
  		c_ap_m1_offsets:missing_value = 65528US, 65529US, 65530US, 65531US, 65532US, 65533US, 65534US, 65535US ;
  		string c_ap_m1_offsets:coordinates = "start_of_scan_time" ;
  		string c_ap_m1_offsets:long_name = "M1 Band FPA Electronics Offsets" ;
  		string c_ap_m1_offsets:source = "APID826:(C_AP_M1_HAM0_DET01-16, C_AP_M1_HAM1_DET01-16)" ;
  	ushort c_ap_m2_offsets(scans, mirror_sides, detectors_750m) ;
  		c_ap_m2_offsets:_FillValue = 65534US ;
  		c_ap_m2_offsets:valid_min = 0US ;
  		c_ap_m2_offsets:valid_max = 65535US ;
  		c_ap_m2_offsets:missing_value = 65528US, 65529US, 65530US, 65531US, 65532US, 65533US, 65534US, 65535US ;
  		string c_ap_m2_offsets:coordinates = "start_of_scan_time" ;
  		string c_ap_m2_offsets:long_name = "M2 Band FPA Electronics Offsets" ;
  		string c_ap_m2_offsets:source = "APID826:(C_AP_M2_HAM0_DET01-16, C_AP_M2_HAM1_DET01-16)" ;
  	ushort c_ap_m3_offsets(scans, mirror_sides, detectors_750m) ;
  		c_ap_m3_offsets:_FillValue = 65534US ;
  		c_ap_m3_offsets:valid_min = 0US ;
  		c_ap_m3_offsets:valid_max = 65535US ;
  		c_ap_m3_offsets:missing_value = 65528US, 65529US, 65530US, 65531US, 65532US, 65533US, 65534US, 65535US ;
  		string c_ap_m3_offsets:coordinates = "start_of_scan_time" ;
  		string c_ap_m3_offsets:long_name = "M3 Band FPA Electronics Offsets" ;
  		string c_ap_m3_offsets:source = "APID826:(C_AP_M3_HAM0_DET01-16, C_AP_M3_HAM1_DET01-16)" ;
  	ushort c_ap_m4_offsets(scans, mirror_sides, detectors_750m) ;
  		c_ap_m4_offsets:_FillValue = 65534US ;
  		c_ap_m4_offsets:valid_min = 0US ;
  		c_ap_m4_offsets:valid_max = 65535US ;
  		c_ap_m4_offsets:missing_value = 65528US, 65529US, 65530US, 65531US, 65532US, 65533US, 65534US, 65535US ;
  		string c_ap_m4_offsets:coordinates = "start_of_scan_time" ;
  		string c_ap_m4_offsets:long_name = "M4 Band FPA Electronics Offsets" ;
  		string c_ap_m4_offsets:source = "APID826:(C_AP_M4_HAM0_DET01-16, C_AP_M4_HAM1_DET01-16)" ;
  	ushort c_ap_m5_offsets(scans, mirror_sides, detectors_750m) ;
  		c_ap_m5_offsets:_FillValue = 65534US ;
  		c_ap_m5_offsets:valid_min = 0US ;
  		c_ap_m5_offsets:valid_max = 65535US ;
  		c_ap_m5_offsets:missing_value = 65528US, 65529US, 65530US, 65531US, 65532US, 65533US, 65534US, 65535US ;
  		string c_ap_m5_offsets:coordinates = "start_of_scan_time" ;
  		string c_ap_m5_offsets:long_name = "M5 Band FPA Electronics Offsets" ;
  		string c_ap_m5_offsets:source = "APID826:(C_AP_M5_HAM0_DET01-16, C_AP_M5_HAM1_DET01-16)" ;
  	ushort c_ap_m6_offsets(scans, mirror_sides, detectors_750m) ;
  		c_ap_m6_offsets:_FillValue = 65534US ;
  		c_ap_m6_offsets:valid_min = 0US ;
  		c_ap_m6_offsets:valid_max = 65535US ;
  		c_ap_m6_offsets:missing_value = 65528US, 65529US, 65530US, 65531US, 65532US, 65533US, 65534US, 65535US ;
  		string c_ap_m6_offsets:coordinates = "start_of_scan_time" ;
  		string c_ap_m6_offsets:long_name = "M6 Band FPA Electronics Offsets" ;
  		string c_ap_m6_offsets:source = "APID826:(C_AP_M6_HAM0_DET01-16, C_AP_M6_HAM1_DET01-16)" ;
  	ushort c_ap_m7_offsets(scans, mirror_sides, detectors_750m) ;
  		c_ap_m7_offsets:_FillValue = 65534US ;
  		c_ap_m7_offsets:valid_min = 0US ;
  		c_ap_m7_offsets:valid_max = 65535US ;
  		c_ap_m7_offsets:missing_value = 65528US, 65529US, 65530US, 65531US, 65532US, 65533US, 65534US, 65535US ;
  		string c_ap_m7_offsets:coordinates = "start_of_scan_time" ;
  		string c_ap_m7_offsets:long_name = "M7 Band FPA Electronics Offsets" ;
  		string c_ap_m7_offsets:source = "APID826:(C_AP_M7_HAM0_DET01-16, C_AP_M7_HAM1_DET01-16)" ;
  	ushort c_ap_m8_offsets(scans, mirror_sides, detectors_750m) ;
  		c_ap_m8_offsets:_FillValue = 65534US ;
  		c_ap_m8_offsets:valid_min = 0US ;
  		c_ap_m8_offsets:valid_max = 65535US ;
  		c_ap_m8_offsets:missing_value = 65528US, 65529US, 65530US, 65531US, 65532US, 65533US, 65534US, 65535US ;
  		string c_ap_m8_offsets:coordinates = "start_of_scan_time" ;
  		string c_ap_m8_offsets:long_name = "M8 Band FPA Electronics Offsets" ;
  		string c_ap_m8_offsets:source = "APID826:(C_AP_M8_HAM0_DET01-16, C_AP_M8_HAM1_DET01-16)" ;
  	ushort c_ap_m9_offsets(scans, mirror_sides, detectors_750m) ;
  		c_ap_m9_offsets:_FillValue = 65534US ;
  		c_ap_m9_offsets:valid_min = 0US ;
  		c_ap_m9_offsets:valid_max = 65535US ;
  		c_ap_m9_offsets:missing_value = 65528US, 65529US, 65530US, 65531US, 65532US, 65533US, 65534US, 65535US ;
  		string c_ap_m9_offsets:coordinates = "start_of_scan_time" ;
  		string c_ap_m9_offsets:long_name = "M9 Band FPA Electronics Offsets" ;
  		string c_ap_m9_offsets:source = "APID826:(C_AP_M9_HAM0_DET01-16, C_AP_M9_HAM1_DET01-16)" ;
  	ushort c_ap_m10_offsets(scans, mirror_sides, detectors_750m) ;
  		c_ap_m10_offsets:_FillValue = 65534US ;
  		c_ap_m10_offsets:valid_min = 0US ;
  		c_ap_m10_offsets:valid_max = 65535US ;
  		c_ap_m10_offsets:missing_value = 65528US, 65529US, 65530US, 65531US, 65532US, 65533US, 65534US, 65535US ;
  		string c_ap_m10_offsets:coordinates = "start_of_scan_time" ;
  		string c_ap_m10_offsets:long_name = "M10 Band FPA Electronics Offsets" ;
  		string c_ap_m10_offsets:source = "APID826:(C_AP_M10_HAM0_DET01-16, C_AP_M10_HAM1_DET01-16)" ;
  	ushort c_ap_m11_offsets(scans, mirror_sides, detectors_750m) ;
  		c_ap_m11_offsets:_FillValue = 65534US ;
  		c_ap_m11_offsets:valid_min = 0US ;
  		c_ap_m11_offsets:valid_max = 65535US ;
  		c_ap_m11_offsets:missing_value = 65528US, 65529US, 65530US, 65531US, 65532US, 65533US, 65534US, 65535US ;
  		string c_ap_m11_offsets:coordinates = "start_of_scan_time" ;
  		string c_ap_m11_offsets:long_name = "M11 Band FPA Electronics Offsets" ;
  		string c_ap_m11_offsets:source = "APID826:(C_AP_M11_HAM0_DET01-16, C_AP_M11_HAM1_DET01-16)" ;
  	ushort c_ap_m12_offsets(scans, mirror_sides, detectors_750m) ;
  		c_ap_m12_offsets:_FillValue = 65534US ;
  		c_ap_m12_offsets:valid_min = 0US ;
  		c_ap_m12_offsets:valid_max = 65535US ;
  		c_ap_m12_offsets:missing_value = 65528US, 65529US, 65530US, 65531US, 65532US, 65533US, 65534US, 65535US ;
  		string c_ap_m12_offsets:coordinates = "start_of_scan_time" ;
  		string c_ap_m12_offsets:long_name = "M12 Band FPA Electronics Offsets" ;
  		string c_ap_m12_offsets:source = "APID826:(C_AP_M12_HAM0_DET01-16, C_AP_M12_HAM1_DET01-16)" ;
  	ushort c_ap_m13_offsets(scans, mirror_sides, detectors_750m) ;
  		c_ap_m13_offsets:_FillValue = 65534US ;
  		c_ap_m13_offsets:valid_min = 0US ;
  		c_ap_m13_offsets:valid_max = 65535US ;
  		c_ap_m13_offsets:missing_value = 65528US, 65529US, 65530US, 65531US, 65532US, 65533US, 65534US, 65535US ;
  		string c_ap_m13_offsets:coordinates = "start_of_scan_time" ;
  		string c_ap_m13_offsets:long_name = "M13 Band FPA Electronics Offsets" ;
  		string c_ap_m13_offsets:source = "APID826:(C_AP_M13_HAM0_DET01-16, C_AP_M13_HAM1_DET01-16)" ;
  	ushort c_ap_m14_offsets(scans, mirror_sides, detectors_750m) ;
  		c_ap_m14_offsets:_FillValue = 65534US ;
  		c_ap_m14_offsets:valid_min = 0US ;
  		c_ap_m14_offsets:valid_max = 65535US ;
  		c_ap_m14_offsets:missing_value = 65528US, 65529US, 65530US, 65531US, 65532US, 65533US, 65534US, 65535US ;
  		string c_ap_m14_offsets:coordinates = "start_of_scan_time" ;
  		string c_ap_m14_offsets:long_name = "M14 Band FPA Electronics Offsets" ;
  		string c_ap_m14_offsets:source = "APID826:(C_AP_M14_HAM0_DET01-16, C_AP_M14_HAM1_DET01-16)" ;
  	ushort c_ap_m15_offsets(scans, mirror_sides, detectors_750m) ;
  		c_ap_m15_offsets:_FillValue = 65534US ;
  		c_ap_m15_offsets:valid_min = 0US ;
  		c_ap_m15_offsets:valid_max = 65535US ;
  		c_ap_m15_offsets:missing_value = 65528US, 65529US, 65530US, 65531US, 65532US, 65533US, 65534US, 65535US ;
  		string c_ap_m15_offsets:coordinates = "start_of_scan_time" ;
  		string c_ap_m15_offsets:long_name = "M15 Band FPA Electronics Offsets" ;
  		string c_ap_m15_offsets:source = "APID826:(C_AP_M15_HAM0_DET01-16, C_AP_M15_HAM1_DET01-16)" ;
  	ushort c_ap_m16a_offsets(scans, mirror_sides, detectors_750m) ;
  		c_ap_m16a_offsets:_FillValue = 65534US ;
  		c_ap_m16a_offsets:valid_min = 0US ;
  		c_ap_m16a_offsets:valid_max = 65535US ;
  		c_ap_m16a_offsets:missing_value = 65528US, 65529US, 65530US, 65531US, 65532US, 65533US, 65534US, 65535US ;
  		string c_ap_m16a_offsets:coordinates = "start_of_scan_time" ;
  		string c_ap_m16a_offsets:long_name = "M16a Band FPA Electronics Offsets" ;
  		string c_ap_m16a_offsets:source = "APID826:(C_AP_M16A_HAM0_DET01-16, C_AP_M16A_HAM1_DET01-16)" ;
  	ushort c_ap_m16b_offsets(scans, mirror_sides, detectors_750m) ;
  		c_ap_m16b_offsets:_FillValue = 65534US ;
  		c_ap_m16b_offsets:valid_min = 0US ;
  		c_ap_m16b_offsets:valid_max = 65535US ;
  		c_ap_m16b_offsets:missing_value = 65528US, 65529US, 65530US, 65531US, 65532US, 65533US, 65534US, 65535US ;
  		string c_ap_m16b_offsets:coordinates = "start_of_scan_time" ;
  		string c_ap_m16b_offsets:long_name = "M16b Band FPA Electronics Offsets" ;
  		string c_ap_m16b_offsets:source = "APID826:(C_AP_M16B_HAM0_DET01-16, C_AP_M16B_HAM1_DET01-16)" ;
  	ushort c_ap_i1_offsets(scans, mirror_sides, detectors_375m) ;
  		c_ap_i1_offsets:_FillValue = 65534US ;
  		c_ap_i1_offsets:valid_min = 0US ;
  		c_ap_i1_offsets:valid_max = 65535US ;
  		c_ap_i1_offsets:missing_value = 65528US, 65529US, 65530US, 65531US, 65532US, 65533US, 65534US, 65535US ;
  		string c_ap_i1_offsets:coordinates = "start_of_scan_time" ;
  		string c_ap_i1_offsets:long_name = "I1 Band FPA Electronics Offsets" ;
  		string c_ap_i1_offsets:source = "APID826:(C_AP_I1E_HAM0_DET01-16, C_AP_I1O_HAM0_DET01-16, C_AP_I1E_HAM1_DET01-16, C_AP_I1O_HAM1_DET01-16)" ;
  	ushort c_ap_i2_offsets(scans, mirror_sides, detectors_375m) ;
  		c_ap_i2_offsets:_FillValue = 65534US ;
  		c_ap_i2_offsets:valid_min = 0US ;
  		c_ap_i2_offsets:valid_max = 65535US ;
  		c_ap_i2_offsets:missing_value = 65528US, 65529US, 65530US, 65531US, 65532US, 65533US, 65534US, 65535US ;
  		string c_ap_i2_offsets:coordinates = "start_of_scan_time" ;
  		string c_ap_i2_offsets:long_name = "I2 Band FPA Electronics Offsets" ;
  		string c_ap_i2_offsets:source = "APID826:(C_AP_I2E_HAM0_DET01-16, C_AP_I2O_HAM0_DET01-16, C_AP_I2E_HAM1_DET01-16, C_AP_I2O_HAM1_DET01-16)" ;
  	ushort c_ap_i3_offsets(scans, mirror_sides, detectors_375m) ;
  		c_ap_i3_offsets:_FillValue = 65534US ;
  		c_ap_i3_offsets:valid_min = 0US ;
  		c_ap_i3_offsets:valid_max = 65535US ;
  		c_ap_i3_offsets:missing_value = 65528US, 65529US, 65530US, 65531US, 65532US, 65533US, 65534US, 65535US ;
  		string c_ap_i3_offsets:coordinates = "start_of_scan_time" ;
  		string c_ap_i3_offsets:long_name = "I3 Band FPA Electronics Offsets" ;
  		string c_ap_i3_offsets:source = "APID826:(C_AP_I3E_HAM0_DET01-16, C_AP_I3O_HAM0_DET01-16, C_AP_I3E_HAM1_DET01-16, C_AP_I3O_HAM1_DET01-16)" ;
  	ushort c_ap_i4_offsets(scans, mirror_sides, detectors_375m) ;
  		c_ap_i4_offsets:_FillValue = 65534US ;
  		c_ap_i4_offsets:valid_min = 0US ;
  		c_ap_i4_offsets:valid_max = 65535US ;
  		c_ap_i4_offsets:missing_value = 65528US, 65529US, 65530US, 65531US, 65532US, 65533US, 65534US, 65535US ;
  		string c_ap_i4_offsets:coordinates = "start_of_scan_time" ;
  		string c_ap_i4_offsets:long_name = "I4 Band FPA Electronics Offsets" ;
  		string c_ap_i4_offsets:source = "APID826:(C_AP_I4E_HAM0_DET01-16, C_AP_I4O_HAM0_DET01-16, C_AP_I4E_HAM1_DET01-16, C_AP_I4O_HAM1_DET01-16)" ;
  	ushort c_ap_i5_offsets(scans, mirror_sides, detectors_375m) ;
  		c_ap_i5_offsets:_FillValue = 65534US ;
  		c_ap_i5_offsets:valid_min = 0US ;
  		c_ap_i5_offsets:valid_max = 65535US ;
  		c_ap_i5_offsets:missing_value = 65528US, 65529US, 65530US, 65531US, 65532US, 65533US, 65534US, 65535US ;
  		string c_ap_i5_offsets:coordinates = "start_of_scan_time" ;
  		string c_ap_i5_offsets:long_name = "I5 Band FPA Electronics Offsets" ;
  		string c_ap_i5_offsets:source = "APID826:(C_AP_I5E_HAM0_DET01-16, C_AP_I5O_HAM0_DET01-16, C_AP_I5E_HAM1_DET01-16, C_AP_I5O_HAM1_DET01-16)" ;
  	ubyte s_cp_events_table(scans, events, event_bytes) ;
  		s_cp_events_table:_FillValue = 254UB ;
  		s_cp_events_table:valid_min = 0UB ;
  		s_cp_events_table:valid_max = 255UB ;
  		s_cp_events_table:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string s_cp_events_table:coordinates = "start_of_scan_time" ;
  		string s_cp_events_table:long_name = "Event Table Dump" ;
  		string s_cp_events_table:source = "APID826:S_CP_EVENTS_TABLE" ;
  	short ev_ap_p30_vispin(scans) ;
  		ev_ap_p30_vispin:_FillValue = -998s ;
  		ev_ap_p30_vispin:valid_min = -8192s ;
  		ev_ap_p30_vispin:valid_max = 8191s ;
  		ev_ap_p30_vispin:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string ev_ap_p30_vispin:coordinates = "start_of_scan_time" ;
  		string ev_ap_p30_vispin:long_name = "Visible/NIR P30_VISPIN Backplane Source Voltage" ;
  		string ev_ap_p30_vispin:source = "APID826:EV_AP_P30_VISPIN" ;
  	short v_ap_lwir_adj_bias_1v(scans) ;
  		v_ap_lwir_adj_bias_1v:_FillValue = -998s ;
  		v_ap_lwir_adj_bias_1v:valid_min = -8192s ;
  		v_ap_lwir_adj_bias_1v:valid_max = 8191s ;
  		v_ap_lwir_adj_bias_1v:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string v_ap_lwir_adj_bias_1v:coordinates = "start_of_scan_time" ;
  		string v_ap_lwir_adj_bias_1v:long_name = "LW-IR Adjust 1V Bias Voltage" ;
  		string v_ap_lwir_adj_bias_1v:source = "APID826:V_AP_LWIR_ADJ_BIAS_1V" ;
  	short v_ap_lwir_adj_bias_2v(scans) ;
  		v_ap_lwir_adj_bias_2v:_FillValue = -998s ;
  		v_ap_lwir_adj_bias_2v:valid_min = -8192s ;
  		v_ap_lwir_adj_bias_2v:valid_max = 8191s ;
  		v_ap_lwir_adj_bias_2v:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string v_ap_lwir_adj_bias_2v:coordinates = "start_of_scan_time" ;
  		string v_ap_lwir_adj_bias_2v:long_name = "LW-IR Adjust 2V Bias Voltage" ;
  		string v_ap_lwir_adj_bias_2v:source = "APID826:V_AP_LWIR_ADJ_BIAS_2V" ;
  	short v_ap_lw_vdet_com1(scans) ;
  		v_ap_lw_vdet_com1:_FillValue = -998s ;
  		v_ap_lw_vdet_com1:valid_min = -8192s ;
  		v_ap_lw_vdet_com1:valid_max = 8191s ;
  		v_ap_lw_vdet_com1:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string v_ap_lw_vdet_com1:coordinates = "start_of_scan_time" ;
  		string v_ap_lw_vdet_com1:long_name = "LW-IR VDET COM1 Bias Voltage" ;
  		string v_ap_lw_vdet_com1:source = "APID826:V_AP_LW_VDET_COM1" ;
  	short v_ap_lw_vdet_com2(scans) ;
  		v_ap_lw_vdet_com2:_FillValue = -998s ;
  		v_ap_lw_vdet_com2:valid_min = -8192s ;
  		v_ap_lw_vdet_com2:valid_max = 8191s ;
  		v_ap_lw_vdet_com2:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string v_ap_lw_vdet_com2:coordinates = "start_of_scan_time" ;
  		string v_ap_lw_vdet_com2:long_name = "LW-IR VDET COM2 Bias Voltage" ;
  		string v_ap_lw_vdet_com2:source = "APID826:V_AP_LW_VDET_COM2" ;
  	short v_ap_lw_vr_clamp(scans) ;
  		v_ap_lw_vr_clamp:_FillValue = -998s ;
  		v_ap_lw_vr_clamp:valid_min = -8192s ;
  		v_ap_lw_vr_clamp:valid_max = 8191s ;
  		v_ap_lw_vr_clamp:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string v_ap_lw_vr_clamp:coordinates = "start_of_scan_time" ;
  		string v_ap_lw_vr_clamp:long_name = "LW-IR VR Clamp Bias Voltage" ;
  		string v_ap_lw_vr_clamp:source = "APID826:V_AP_LW_VR_CLAMP" ;
  	short v_ap_lw_vi_clamp(scans) ;
  		v_ap_lw_vi_clamp:_FillValue = -998s ;
  		v_ap_lw_vi_clamp:valid_min = -8192s ;
  		v_ap_lw_vi_clamp:valid_max = 8191s ;
  		v_ap_lw_vi_clamp:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string v_ap_lw_vi_clamp:coordinates = "start_of_scan_time" ;
  		string v_ap_lw_vi_clamp:long_name = "LW-IR VI Clamp Bias Voltage" ;
  		string v_ap_lw_vi_clamp:source = "APID826:V_AP_LW_VI_CLAMP" ;
  	short v_ap_lw_vpo(scans) ;
  		v_ap_lw_vpo:_FillValue = -998s ;
  		v_ap_lw_vpo:valid_min = -8192s ;
  		v_ap_lw_vpo:valid_max = 8191s ;
  		v_ap_lw_vpo:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string v_ap_lw_vpo:coordinates = "start_of_scan_time" ;
  		string v_ap_lw_vpo:long_name = "LW-IR VPO Bias Voltage" ;
  		string v_ap_lw_vpo:source = "APID826:V_AP_LW_VPO" ;
  	short v_ap_lw_vna(scans) ;
  		v_ap_lw_vna:_FillValue = -998s ;
  		v_ap_lw_vna:valid_min = -8192s ;
  		v_ap_lw_vna:valid_max = 8191s ;
  		v_ap_lw_vna:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string v_ap_lw_vna:coordinates = "start_of_scan_time" ;
  		string v_ap_lw_vna:long_name = "LW-IR VNA Bias Voltage" ;
  		string v_ap_lw_vna:source = "APID826:V_AP_LW_VNA" ;
  	short v_ap_lw_vnd(scans) ;
  		v_ap_lw_vnd:_FillValue = -998s ;
  		v_ap_lw_vnd:valid_min = -8192s ;
  		v_ap_lw_vnd:valid_max = 8191s ;
  		v_ap_lw_vnd:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string v_ap_lw_vnd:coordinates = "start_of_scan_time" ;
  		string v_ap_lw_vnd:long_name = "LW-IR VND Bias Voltage" ;
  		string v_ap_lw_vnd:source = "APID826:V_AP_LW_VND" ;
  	short v_ap_lw_vn_stat(scans) ;
  		v_ap_lw_vn_stat:_FillValue = -998s ;
  		v_ap_lw_vn_stat:valid_min = -8192s ;
  		v_ap_lw_vn_stat:valid_max = 8191s ;
  		v_ap_lw_vn_stat:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string v_ap_lw_vn_stat:coordinates = "start_of_scan_time" ;
  		string v_ap_lw_vn_stat:long_name = "LW-IR VN Stat Bias Voltage" ;
  		string v_ap_lw_vn_stat:source = "APID826:V_AP_LW_VN_STAT" ;
  	short v_ap_smwir_adj_bias_1v(scans) ;
  		v_ap_smwir_adj_bias_1v:_FillValue = -998s ;
  		v_ap_smwir_adj_bias_1v:valid_min = -8192s ;
  		v_ap_smwir_adj_bias_1v:valid_max = 8191s ;
  		v_ap_smwir_adj_bias_1v:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string v_ap_smwir_adj_bias_1v:coordinates = "start_of_scan_time" ;
  		string v_ap_smwir_adj_bias_1v:long_name = "SW/MW-IR Adjust 1V Bias Voltage" ;
  		string v_ap_smwir_adj_bias_1v:source = "APID826:V_AP_SMWIR_ADJ_BIAS_1V" ;
  	short v_ap_smwir_adj_bias_2v(scans) ;
  		v_ap_smwir_adj_bias_2v:_FillValue = -998s ;
  		v_ap_smwir_adj_bias_2v:valid_min = -8192s ;
  		v_ap_smwir_adj_bias_2v:valid_max = 8191s ;
  		v_ap_smwir_adj_bias_2v:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string v_ap_smwir_adj_bias_2v:coordinates = "start_of_scan_time" ;
  		string v_ap_smwir_adj_bias_2v:long_name = "SW/MW-IR Adjust 2V Bias Voltage" ;
  		string v_ap_smwir_adj_bias_2v:source = "APID826:V_AP_SMWIR_ADJ_BIAS_2V" ;
  	short v_ap_sm_vnrst(scans) ;
  		v_ap_sm_vnrst:_FillValue = -998s ;
  		v_ap_sm_vnrst:valid_min = -8192s ;
  		v_ap_sm_vnrst:valid_max = 8191s ;
  		v_ap_sm_vnrst:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string v_ap_sm_vnrst:coordinates = "start_of_scan_time" ;
  		string v_ap_sm_vnrst:long_name = "SW/MW-IR VNRST Bias Voltage" ;
  		string v_ap_sm_vnrst:source = "APID826:V_AP_SM_VNRST" ;
  	short v_ap_sm_dgain_sw_vref(scans) ;
  		v_ap_sm_dgain_sw_vref:_FillValue = -998s ;
  		v_ap_sm_dgain_sw_vref:valid_min = -8192s ;
  		v_ap_sm_dgain_sw_vref:valid_max = 8191s ;
  		v_ap_sm_dgain_sw_vref:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string v_ap_sm_dgain_sw_vref:coordinates = "start_of_scan_time" ;
  		string v_ap_sm_dgain_sw_vref:long_name = "SW/MW-IR Dual Gain Transition Bias Voltage" ;
  		string v_ap_sm_dgain_sw_vref:source = "APID826:V_AP_SM_DGAIN_SW_VREF" ;
  	short v_ap_sm_vr_clamp(scans) ;
  		v_ap_sm_vr_clamp:_FillValue = -998s ;
  		v_ap_sm_vr_clamp:valid_min = -8192s ;
  		v_ap_sm_vr_clamp:valid_max = 8191s ;
  		v_ap_sm_vr_clamp:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string v_ap_sm_vr_clamp:coordinates = "start_of_scan_time" ;
  		string v_ap_sm_vr_clamp:long_name = "SW/MW-IR VR Clamp Bias Voltage" ;
  		string v_ap_sm_vr_clamp:source = "APID826:V_AP_SM_VR_CLAMP" ;
  	short v_ap_sm_vi_clamp(scans) ;
  		v_ap_sm_vi_clamp:_FillValue = -998s ;
  		v_ap_sm_vi_clamp:valid_min = -8192s ;
  		v_ap_sm_vi_clamp:valid_max = 8191s ;
  		v_ap_sm_vi_clamp:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string v_ap_sm_vi_clamp:coordinates = "start_of_scan_time" ;
  		string v_ap_sm_vi_clamp:long_name = "SW/MW-IR VI Clamp Bias Voltage" ;
  		string v_ap_sm_vi_clamp:source = "APID826:V_AP_SM_VI_CLAMP" ;
  	short v_ap_sm_vpo(scans) ;
  		v_ap_sm_vpo:_FillValue = -998s ;
  		v_ap_sm_vpo:valid_min = -8192s ;
  		v_ap_sm_vpo:valid_max = 8191s ;
  		v_ap_sm_vpo:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string v_ap_sm_vpo:coordinates = "start_of_scan_time" ;
  		string v_ap_sm_vpo:long_name = "SW/MW-IR VPO Bias Voltage" ;
  		string v_ap_sm_vpo:source = "APID826:V_AP_SM_VPO" ;
  	short v_ap_sm_vna(scans) ;
  		v_ap_sm_vna:_FillValue = -998s ;
  		v_ap_sm_vna:valid_min = -8192s ;
  		v_ap_sm_vna:valid_max = 8191s ;
  		v_ap_sm_vna:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string v_ap_sm_vna:coordinates = "start_of_scan_time" ;
  		string v_ap_sm_vna:long_name = "SW/MW-IR VNA Bias Voltage" ;
  		string v_ap_sm_vna:source = "APID826:V_AP_SM_VNA" ;
  	short v_ap_sm_vnd(scans) ;
  		v_ap_sm_vnd:_FillValue = -998s ;
  		v_ap_sm_vnd:valid_min = -8192s ;
  		v_ap_sm_vnd:valid_max = 8191s ;
  		v_ap_sm_vnd:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string v_ap_sm_vnd:coordinates = "start_of_scan_time" ;
  		string v_ap_sm_vnd:long_name = "SW/MW-IR VND Bias Voltage" ;
  		string v_ap_sm_vnd:source = "APID826:V_AP_SM_VND" ;
  	short v_ap_sm_vn_stat(scans) ;
  		v_ap_sm_vn_stat:_FillValue = -998s ;
  		v_ap_sm_vn_stat:valid_min = -8192s ;
  		v_ap_sm_vn_stat:valid_max = 8191s ;
  		v_ap_sm_vn_stat:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string v_ap_sm_vn_stat:coordinates = "start_of_scan_time" ;
  		string v_ap_sm_vn_stat:long_name = "SW/MW-IR VN Stat Bias Voltage" ;
  		string v_ap_sm_vn_stat:source = "APID826:V_AP_SM_VN_STAT" ;
  	short v_ap_visnir_adj_bias_1v(scans) ;
  		v_ap_visnir_adj_bias_1v:_FillValue = -998s ;
  		v_ap_visnir_adj_bias_1v:valid_min = -8192s ;
  		v_ap_visnir_adj_bias_1v:valid_max = 8191s ;
  		v_ap_visnir_adj_bias_1v:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string v_ap_visnir_adj_bias_1v:coordinates = "start_of_scan_time" ;
  		string v_ap_visnir_adj_bias_1v:long_name = "Visible/NIR Adjust 1V Bias Voltage" ;
  		string v_ap_visnir_adj_bias_1v:source = "APID826:V_AP_VISNIR_ADJ_BIAS_1V" ;
  	short ev_ap_vn_dgain_sw_vref(scans) ;
  		ev_ap_vn_dgain_sw_vref:_FillValue = -998s ;
  		ev_ap_vn_dgain_sw_vref:valid_min = -8192s ;
  		ev_ap_vn_dgain_sw_vref:valid_max = 8191s ;
  		ev_ap_vn_dgain_sw_vref:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string ev_ap_vn_dgain_sw_vref:coordinates = "start_of_scan_time" ;
  		string ev_ap_vn_dgain_sw_vref:long_name = "Visible/NIR Dual Gain Transition Bias Voltage" ;
  		string ev_ap_vn_dgain_sw_vref:source = "APID826:EV_AP_VN_DGAIN_SW_VREF" ;
  	short v_ap_vn_vdet_com1(scans) ;
  		v_ap_vn_vdet_com1:_FillValue = -998s ;
  		v_ap_vn_vdet_com1:valid_min = -8192s ;
  		v_ap_vn_vdet_com1:valid_max = 8191s ;
  		v_ap_vn_vdet_com1:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string v_ap_vn_vdet_com1:coordinates = "start_of_scan_time" ;
  		string v_ap_vn_vdet_com1:long_name = "Visible/NIR VDET COM1 Bias Voltage" ;
  		string v_ap_vn_vdet_com1:source = "APID826:V_AP_VN_VDET_COM1" ;
  	short v_ap_vn_vdet_com2(scans) ;
  		v_ap_vn_vdet_com2:_FillValue = -998s ;
  		v_ap_vn_vdet_com2:valid_min = -8192s ;
  		v_ap_vn_vdet_com2:valid_max = 8191s ;
  		v_ap_vn_vdet_com2:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string v_ap_vn_vdet_com2:coordinates = "start_of_scan_time" ;
  		string v_ap_vn_vdet_com2:long_name = "Visible/NIR VDET COM2 Bias Voltage" ;
  		string v_ap_vn_vdet_com2:source = "APID826:V_AP_VN_VDET_COM2" ;
  	short v_ap_vn_vr_clamp(scans) ;
  		v_ap_vn_vr_clamp:_FillValue = -998s ;
  		v_ap_vn_vr_clamp:valid_min = -8192s ;
  		v_ap_vn_vr_clamp:valid_max = 8191s ;
  		v_ap_vn_vr_clamp:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string v_ap_vn_vr_clamp:coordinates = "start_of_scan_time" ;
  		string v_ap_vn_vr_clamp:long_name = "Visible/NIR VR Clamp Bias Voltage" ;
  		string v_ap_vn_vr_clamp:source = "APID826:V_AP_VN_VR_CLAMP" ;
  	short v_ap_vn_vi_clamp(scans) ;
  		v_ap_vn_vi_clamp:_FillValue = -998s ;
  		v_ap_vn_vi_clamp:valid_min = -8192s ;
  		v_ap_vn_vi_clamp:valid_max = 8191s ;
  		v_ap_vn_vi_clamp:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string v_ap_vn_vi_clamp:coordinates = "start_of_scan_time" ;
  		string v_ap_vn_vi_clamp:long_name = "Visible/NIR VI Clamp Bias Voltage" ;
  		string v_ap_vn_vi_clamp:source = "APID826:V_AP_VN_VI_CLAMP" ;
  	short v_ap_vn_vpo(scans) ;
  		v_ap_vn_vpo:_FillValue = -998s ;
  		v_ap_vn_vpo:valid_min = -8192s ;
  		v_ap_vn_vpo:valid_max = 8191s ;
  		v_ap_vn_vpo:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string v_ap_vn_vpo:coordinates = "start_of_scan_time" ;
  		string v_ap_vn_vpo:long_name = "Visible/NIR VPO Bias Voltage" ;
  		string v_ap_vn_vpo:source = "APID826:V_AP_VN_VPO" ;
  	short v_ap_vn_vna(scans) ;
  		v_ap_vn_vna:_FillValue = -998s ;
  		v_ap_vn_vna:valid_min = -8192s ;
  		v_ap_vn_vna:valid_max = 8191s ;
  		v_ap_vn_vna:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string v_ap_vn_vna:coordinates = "start_of_scan_time" ;
  		string v_ap_vn_vna:long_name = "Visible/NIR VNA Bias Voltage" ;
  		string v_ap_vn_vna:source = "APID826:V_AP_VN_VNA" ;
  	short v_ap_vn_vnd(scans) ;
  		v_ap_vn_vnd:_FillValue = -998s ;
  		v_ap_vn_vnd:valid_min = -8192s ;
  		v_ap_vn_vnd:valid_max = 8191s ;
  		v_ap_vn_vnd:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string v_ap_vn_vnd:coordinates = "start_of_scan_time" ;
  		string v_ap_vn_vnd:long_name = "Visible/NIR VND Bias Voltage" ;
  		string v_ap_vn_vnd:source = "APID826:V_AP_VN_VND" ;
  	short v_ap_vn_vn_stat(scans) ;
  		v_ap_vn_vn_stat:_FillValue = -998s ;
  		v_ap_vn_vn_stat:valid_min = -8192s ;
  		v_ap_vn_vn_stat:valid_max = 8191s ;
  		v_ap_vn_vn_stat:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string v_ap_vn_vn_stat:coordinates = "start_of_scan_time" ;
  		string v_ap_vn_vn_stat:long_name = "Visible/NIR VN Stat Bias Voltage" ;
  		string v_ap_vn_vn_stat:source = "APID826:V_AP_VN_VN_STAT" ;
  	ushort ec_ap_lw_selftest_vb(scans) ;
  		ec_ap_lw_selftest_vb:_FillValue = 65534US ;
  		ec_ap_lw_selftest_vb:valid_min = 0US ;
  		ec_ap_lw_selftest_vb:valid_max = 4095US ;
  		ec_ap_lw_selftest_vb:missing_value = 65528US, 65529US, 65530US, 65531US, 65532US, 65533US, 65534US, 65535US ;
  		string ec_ap_lw_selftest_vb:coordinates = "start_of_scan_time" ;
  		string ec_ap_lw_selftest_vb:long_name = "LW-IR Self-test Commanded Vbase Voltage" ;
  		string ec_ap_lw_selftest_vb:source = "APID826:EC_AP_LW_SELFTEST_VB" ;
  	ushort ec_ap_lw_selftest_vs_cm(scans) ;
  		ec_ap_lw_selftest_vs_cm:_FillValue = 65534US ;
  		ec_ap_lw_selftest_vs_cm:valid_min = 0US ;
  		ec_ap_lw_selftest_vs_cm:valid_max = 4095US ;
  		ec_ap_lw_selftest_vs_cm:missing_value = 65528US, 65529US, 65530US, 65531US, 65532US, 65533US, 65534US, 65535US ;
  		string ec_ap_lw_selftest_vs_cm:coordinates = "start_of_scan_time" ;
  		string ec_ap_lw_selftest_vs_cm:long_name = "LW-IR Self-test Commanded Vstep Voltage" ;
  		string ec_ap_lw_selftest_vs_cm:source = "APID826:EC_AP_LW_SELFTEST_VS_CM" ;
  	short ev_ap_lw_selftest_vs_tl(scans) ;
  		ev_ap_lw_selftest_vs_tl:_FillValue = -998s ;
  		ev_ap_lw_selftest_vs_tl:valid_min = -8192s ;
  		ev_ap_lw_selftest_vs_tl:valid_max = 8191s ;
  		ev_ap_lw_selftest_vs_tl:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string ev_ap_lw_selftest_vs_tl:coordinates = "start_of_scan_time" ;
  		string ev_ap_lw_selftest_vs_tl:long_name = "LW-IR Self-test Vstep Voltage" ;
  		string ev_ap_lw_selftest_vs_tl:source = "APID826:EV_AP_LW_SELFTEST_VS_TL" ;
  	short ev_ap_lw_vab_adj(scans) ;
  		ev_ap_lw_vab_adj:_FillValue = -998s ;
  		ev_ap_lw_vab_adj:valid_min = -8192s ;
  		ev_ap_lw_vab_adj:valid_max = 8191s ;
  		ev_ap_lw_vab_adj:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string ev_ap_lw_vab_adj:coordinates = "start_of_scan_time" ;
  		string ev_ap_lw_vab_adj:long_name = "LW-IR FPA Variable Detector Bias Voltage" ;
  		string ev_ap_lw_vab_adj:source = "APID826:EV_AP_LW_VAB_ADJ" ;
  	short ev_ap_lw_vdet_adj(scans) ;
  		ev_ap_lw_vdet_adj:_FillValue = -998s ;
  		ev_ap_lw_vdet_adj:valid_min = -8192s ;
  		ev_ap_lw_vdet_adj:valid_max = 8191s ;
  		ev_ap_lw_vdet_adj:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string ev_ap_lw_vdet_adj:coordinates = "start_of_scan_time" ;
  		string ev_ap_lw_vdet_adj:long_name = "LW-IR FPA Fixed Detector Bias Voltage" ;
  		string ev_ap_lw_vdet_adj:source = "APID826:EV_AP_LW_VDET_ADJ" ;
  	ushort ec_ap_sm_selftest_vb(scans) ;
  		ec_ap_sm_selftest_vb:_FillValue = 65534US ;
  		ec_ap_sm_selftest_vb:valid_min = 0US ;
  		ec_ap_sm_selftest_vb:valid_max = 4095US ;
  		ec_ap_sm_selftest_vb:missing_value = 65528US, 65529US, 65530US, 65531US, 65532US, 65533US, 65534US, 65535US ;
  		string ec_ap_sm_selftest_vb:coordinates = "start_of_scan_time" ;
  		string ec_ap_sm_selftest_vb:long_name = "SW/MW-IR Self-test Commanded Vbase Voltage" ;
  		string ec_ap_sm_selftest_vb:source = "APID826:EC_AP_SM_SELFTEST_VB" ;
  	ushort ec_ap_sm_selftest_vs_cm(scans) ;
  		ec_ap_sm_selftest_vs_cm:_FillValue = 65534US ;
  		ec_ap_sm_selftest_vs_cm:valid_min = 0US ;
  		ec_ap_sm_selftest_vs_cm:valid_max = 4095US ;
  		ec_ap_sm_selftest_vs_cm:missing_value = 65528US, 65529US, 65530US, 65531US, 65532US, 65533US, 65534US, 65535US ;
  		string ec_ap_sm_selftest_vs_cm:coordinates = "start_of_scan_time" ;
  		string ec_ap_sm_selftest_vs_cm:long_name = "SW/MW-IR Self-test Commanded Vstep Voltage" ;
  		string ec_ap_sm_selftest_vs_cm:source = "APID826:EC_AP_SM_SELFTEST_VS_CM" ;
  	short ev_ap_sm_selftest_vs_tl(scans) ;
  		ev_ap_sm_selftest_vs_tl:_FillValue = -998s ;
  		ev_ap_sm_selftest_vs_tl:valid_min = -8192s ;
  		ev_ap_sm_selftest_vs_tl:valid_max = 8191s ;
  		ev_ap_sm_selftest_vs_tl:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string ev_ap_sm_selftest_vs_tl:coordinates = "start_of_scan_time" ;
  		string ev_ap_sm_selftest_vs_tl:long_name = "SW/MW-IR Self-test Vstep Voltage" ;
  		string ev_ap_sm_selftest_vs_tl:source = "APID826:EV_AP_SM_SELFTEST_VS_TL" ;
  	short ev_ap_sm_vab_adj(scans) ;
  		ev_ap_sm_vab_adj:_FillValue = -998s ;
  		ev_ap_sm_vab_adj:valid_min = -8192s ;
  		ev_ap_sm_vab_adj:valid_max = 8191s ;
  		ev_ap_sm_vab_adj:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string ev_ap_sm_vab_adj:coordinates = "start_of_scan_time" ;
  		string ev_ap_sm_vab_adj:long_name = "SW/MW-IR FPA Variable Detector Bias Voltage" ;
  		string ev_ap_sm_vab_adj:source = "APID826:EV_AP_SM_VAB_ADJ" ;
  	short ev_ap_sm_dgain_sw_vref(scans) ;
  		ev_ap_sm_dgain_sw_vref:_FillValue = -998s ;
  		ev_ap_sm_dgain_sw_vref:valid_min = -8192s ;
  		ev_ap_sm_dgain_sw_vref:valid_max = 8191s ;
  		ev_ap_sm_dgain_sw_vref:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string ev_ap_sm_dgain_sw_vref:coordinates = "start_of_scan_time" ;
  		string ev_ap_sm_dgain_sw_vref:long_name = "SW/MW-IR Dual Gain Transition Bias Voltage (copy)" ;
  		string ev_ap_sm_dgain_sw_vref:source = "APID826:EV_AP_SM_DGAIN_SW_VREF" ;
  	ushort ec_ap_vn_selftest_vb(scans) ;
  		ec_ap_vn_selftest_vb:_FillValue = 65534US ;
  		ec_ap_vn_selftest_vb:valid_min = 0US ;
  		ec_ap_vn_selftest_vb:valid_max = 4095US ;
  		ec_ap_vn_selftest_vb:missing_value = 65528US, 65529US, 65530US, 65531US, 65532US, 65533US, 65534US, 65535US ;
  		string ec_ap_vn_selftest_vb:coordinates = "start_of_scan_time" ;
  		string ec_ap_vn_selftest_vb:long_name = "Visible/NIR Self-test Commanded Vbase Voltage" ;
  		string ec_ap_vn_selftest_vb:source = "APID826:EC_AP_VN_SELFTEST_VB" ;
  	ushort ec_ap_vn_selftest_vs_cm(scans) ;
  		ec_ap_vn_selftest_vs_cm:_FillValue = 65534US ;
  		ec_ap_vn_selftest_vs_cm:valid_min = 0US ;
  		ec_ap_vn_selftest_vs_cm:valid_max = 4095US ;
  		ec_ap_vn_selftest_vs_cm:missing_value = 65528US, 65529US, 65530US, 65531US, 65532US, 65533US, 65534US, 65535US ;
  		string ec_ap_vn_selftest_vs_cm:coordinates = "start_of_scan_time" ;
  		string ec_ap_vn_selftest_vs_cm:long_name = "Visible/NIR Self-test Commanded Vstep Voltage" ;
  		string ec_ap_vn_selftest_vs_cm:source = "APID826:EC_AP_VN_SELFTEST_VS_CM" ;
  	short ev_ap_vn_selftest_vs_tl(scans) ;
  		ev_ap_vn_selftest_vs_tl:_FillValue = -998s ;
  		ev_ap_vn_selftest_vs_tl:valid_min = -8192s ;
  		ev_ap_vn_selftest_vs_tl:valid_max = 8191s ;
  		ev_ap_vn_selftest_vs_tl:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string ev_ap_vn_selftest_vs_tl:coordinates = "start_of_scan_time" ;
  		string ev_ap_vn_selftest_vs_tl:long_name = "Visible/NIR Self-test Vstep Voltage" ;
  		string ev_ap_vn_selftest_vs_tl:source = "APID826:EV_AP_VN_SELFTEST_VS_TL" ;
  	short ev_ap_vn_vab_adj(scans) ;
  		ev_ap_vn_vab_adj:_FillValue = -998s ;
  		ev_ap_vn_vab_adj:valid_min = -8192s ;
  		ev_ap_vn_vab_adj:valid_max = 8191s ;
  		ev_ap_vn_vab_adj:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string ev_ap_vn_vab_adj:coordinates = "start_of_scan_time" ;
  		string ev_ap_vn_vab_adj:long_name = "Visible/NIR FPA Variable Detector Bias Voltage" ;
  		string ev_ap_vn_vab_adj:source = "APID826:EV_AP_VN_VAB_ADJ" ;
  	short etp_bb_temps(scans, bb_thermistors) ;
  		etp_bb_temps:_FillValue = -998s ;
  		etp_bb_temps:valid_min = -8192s ;
  		etp_bb_temps:valid_max = 8191s ;
  		etp_bb_temps:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string etp_bb_temps:coordinates = "start_of_scan_time" ;
  		string etp_bb_temps:long_name = "Blackbody Temperatures (Thermistors 1-6)" ;
  		string etp_bb_temps:source = "APID826:(ETP_BB_1, ETP_BB_2, ETP_BB_3, ETP_BB_4, ETP_BB_5, ETP_BB_6)" ;
  	short etp_se_ham_mirr_t1(scans) ;
  		etp_se_ham_mirr_t1:_FillValue = -998s ;
  		etp_se_ham_mirr_t1:valid_min = -8192s ;
  		etp_se_ham_mirr_t1:valid_max = 8191s ;
  		etp_se_ham_mirr_t1:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string etp_se_ham_mirr_t1:coordinates = "start_of_scan_time" ;
  		string etp_se_ham_mirr_t1:long_name = "Half-Angle Mirror T2 Precision Thermistor 07, Radiatively coupled (used in Radiometry Model)" ;
  		string etp_se_ham_mirr_t1:source = "APID826:ETP_SE_HAM_MIRR_T1" ;
  	short etp_se_ham_mirr_t2(scans) ;
  		etp_se_ham_mirr_t2:_FillValue = -998s ;
  		etp_se_ham_mirr_t2:valid_min = -8192s ;
  		etp_se_ham_mirr_t2:valid_max = 8191s ;
  		etp_se_ham_mirr_t2:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string etp_se_ham_mirr_t2:coordinates = "start_of_scan_time" ;
  		string etp_se_ham_mirr_t2:long_name = "Half-Angle Mirror T2 Precision Thermistor 08, Radiatively coupled (used in Radiometry Model)" ;
  		string etp_se_ham_mirr_t2:source = "APID826:ETP_SE_HAM_MIRR_T2" ;
  	short etp_hm_cr_cs_prt(scans) ;
  		etp_hm_cr_cs_prt:_FillValue = -998s ;
  		etp_hm_cr_cs_prt:valid_min = -8192s ;
  		etp_hm_cr_cs_prt:valid_max = 8191s ;
  		etp_hm_cr_cs_prt:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string etp_hm_cr_cs_prt:coordinates = "start_of_scan_time" ;
  		string etp_hm_cr_cs_prt:long_name = "CR Cold Stage PRT Temperature" ;
  		string etp_hm_cr_cs_prt:source = "APID826:ETA_HM_CR_CS_PRT" ;
  	short etp_hm_cr_is_prt(scans) ;
  		etp_hm_cr_is_prt:_FillValue = -998s ;
  		etp_hm_cr_is_prt:valid_min = -8192s ;
  		etp_hm_cr_is_prt:valid_max = 8191s ;
  		etp_hm_cr_is_prt:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string etp_hm_cr_is_prt:coordinates = "start_of_scan_time" ;
  		string etp_hm_cr_is_prt:long_name = "CR Intermediate Stage PRT Temperature" ;
  		string etp_hm_cr_is_prt:source = "APID826:ETA_HM_CR_IS_PRT" ;
  	short etp_hm_cr_os_prt(scans) ;
  		etp_hm_cr_os_prt:_FillValue = -998s ;
  		etp_hm_cr_os_prt:valid_min = -8192s ;
  		etp_hm_cr_os_prt:valid_max = 8191s ;
  		etp_hm_cr_os_prt:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string etp_hm_cr_os_prt:coordinates = "start_of_scan_time" ;
  		string etp_hm_cr_os_prt:long_name = "CR Outer Stage PRT Temperature" ;
  		string etp_hm_cr_os_prt:source = "APID826:ETA_HM_CR_OS_PRT" ;
  	short ec_ap_vn_vref_inhibit(scans) ;
  		ec_ap_vn_vref_inhibit:_FillValue = -998s ;
  		ec_ap_vn_vref_inhibit:valid_min = -2048s ;
  		ec_ap_vn_vref_inhibit:valid_max = 2047s ;
  		ec_ap_vn_vref_inhibit:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string ec_ap_vn_vref_inhibit:coordinates = "start_of_scan_time" ;
  		string ec_ap_vn_vref_inhibit:long_name = "Visible/NIR Reference Voltage Inhibit Commanded Voltage" ;
  		string ec_ap_vn_vref_inhibit:source = "APID826:EC_AP_VN_VREF_INHIBIT" ;
  	short etp_hm_ham_db_op_htr_a(scans) ;
  		etp_hm_ham_db_op_htr_a:_FillValue = -998s ;
  		etp_hm_ham_db_op_htr_a:valid_min = -8192s ;
  		etp_hm_ham_db_op_htr_a:valid_max = 8191s ;
  		etp_hm_ham_db_op_htr_a:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string etp_hm_ham_db_op_htr_a:coordinates = "start_of_scan_time" ;
  		string etp_hm_ham_db_op_htr_a:long_name = "Half-Angle Mirror DB Bearing Operational Heater A Temperature (Thermistor 17)" ;
  		string etp_hm_ham_db_op_htr_a:source = "APID826:ETP_HM_HAM_DB_OP_HTR_A" ;
  	short etp_hm_ham_db_op_htr_b(scans) ;
  		etp_hm_ham_db_op_htr_b:_FillValue = -998s ;
  		etp_hm_ham_db_op_htr_b:valid_min = -8192s ;
  		etp_hm_ham_db_op_htr_b:valid_max = 8191s ;
  		etp_hm_ham_db_op_htr_b:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string etp_hm_ham_db_op_htr_b:coordinates = "start_of_scan_time" ;
  		string etp_hm_ham_db_op_htr_b:long_name = "Half-Angle Mirror DB Bearing Operational Heater B Temperature (Thermistor 21)" ;
  		string etp_hm_ham_db_op_htr_b:source = "APID826:ETP_HM_HAM_DB_OP_HTR_B" ;
  	short etp_hm_tele_db_op_htr_a(scans) ;
  		etp_hm_tele_db_op_htr_a:_FillValue = -998s ;
  		etp_hm_tele_db_op_htr_a:valid_min = -8192s ;
  		etp_hm_tele_db_op_htr_a:valid_max = 8191s ;
  		etp_hm_tele_db_op_htr_a:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string etp_hm_tele_db_op_htr_a:coordinates = "start_of_scan_time" ;
  		string etp_hm_tele_db_op_htr_a:long_name = "Telescope DB Bearing Operational Heater A Temperature (Thermistor 18)" ;
  		string etp_hm_tele_db_op_htr_a:source = "APID826:ETP_HM_TELE_DB_OP_HTR_A" ;
  	short etp_hm_tele_db_op_htr_b(scans) ;
  		etp_hm_tele_db_op_htr_b:_FillValue = -998s ;
  		etp_hm_tele_db_op_htr_b:valid_min = -8192s ;
  		etp_hm_tele_db_op_htr_b:valid_max = 8191s ;
  		etp_hm_tele_db_op_htr_b:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string etp_hm_tele_db_op_htr_b:coordinates = "start_of_scan_time" ;
  		string etp_hm_tele_db_op_htr_b:long_name = "Telescope DB Bearing Operational Heater A Temperature (Thermistor 23)" ;
  		string etp_hm_tele_db_op_htr_b:source = "APID826:ETP_HM_TELE_DB_OP_HTR_B" ;
  	short etp_mf_ao_blkhd_nx_pz(scans) ;
  		etp_mf_ao_blkhd_nx_pz:_FillValue = -998s ;
  		etp_mf_ao_blkhd_nx_pz:valid_min = -8192s ;
  		etp_mf_ao_blkhd_nx_pz:valid_max = 8191s ;
  		etp_mf_ao_blkhd_nx_pz:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string etp_mf_ao_blkhd_nx_pz:coordinates = "start_of_scan_time" ;
  		string etp_mf_ao_blkhd_nx_pz:long_name = "Aft Optics Bulkhead NX-PZ Temperature (Thermistor 45)" ;
  		string etp_mf_ao_blkhd_nx_pz:source = "APID826:ETP_MF_AO_BLKHD_NX_PZ" ;
  	short etp_mf_ao_blkhd_px_nz(scans) ;
  		etp_mf_ao_blkhd_px_nz:_FillValue = -998s ;
  		etp_mf_ao_blkhd_px_nz:valid_min = -8192s ;
  		etp_mf_ao_blkhd_px_nz:valid_max = 8191s ;
  		etp_mf_ao_blkhd_px_nz:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string etp_mf_ao_blkhd_px_nz:coordinates = "start_of_scan_time" ;
  		string etp_mf_ao_blkhd_px_nz:long_name = "Aft Optics Bulkhead PX-NZ Temperature (Thermistor 44)" ;
  		string etp_mf_ao_blkhd_px_nz:source = "APID826:ETP_MF_AO_BLKHD_PX_NZ" ;
  	short etp_mf_ao_km2_nx(scans) ;
  		etp_mf_ao_km2_nx:_FillValue = -998s ;
  		etp_mf_ao_km2_nx:valid_min = -8192s ;
  		etp_mf_ao_km2_nx:valid_max = 8191s ;
  		etp_mf_ao_km2_nx:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string etp_mf_ao_km2_nx:coordinates = "start_of_scan_time" ;
  		string etp_mf_ao_km2_nx:long_name = "Aft Optics KM2-NX Temperature (Thermistor 88)" ;
  		string etp_mf_ao_km2_nx:source = "APID826:ETP_MF_AO_KM2_NX" ;
  	short etp_mf_ao_km2_ny(scans) ;
  		etp_mf_ao_km2_ny:_FillValue = -998s ;
  		etp_mf_ao_km2_ny:valid_min = -8192s ;
  		etp_mf_ao_km2_ny:valid_max = 8191s ;
  		etp_mf_ao_km2_ny:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string etp_mf_ao_km2_ny:coordinates = "start_of_scan_time" ;
  		string etp_mf_ao_km2_ny:long_name = "Aft Optics KM2-NY Temperature (Thermistor 39)" ;
  		string etp_mf_ao_km2_ny:source = "APID826:ETP_MF_AO_KM2_NY" ;
  	short etp_mf_ao_km3_px(scans) ;
  		etp_mf_ao_km3_px:_FillValue = -998s ;
  		etp_mf_ao_km3_px:valid_min = -8192s ;
  		etp_mf_ao_km3_px:valid_max = 8191s ;
  		etp_mf_ao_km3_px:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string etp_mf_ao_km3_px:coordinates = "start_of_scan_time" ;
  		string etp_mf_ao_km3_px:long_name = "Aft Optics KM3-PX Temperature (Thermistor 40)" ;
  		string etp_mf_ao_km3_px:source = "APID826:ETP_MF_AO_KM3_PX" ;
  	short etp_mf_fold_mir_bkhd_ct(scans) ;
  		etp_mf_fold_mir_bkhd_ct:_FillValue = -998s ;
  		etp_mf_fold_mir_bkhd_ct:valid_min = -8192s ;
  		etp_mf_fold_mir_bkhd_ct:valid_max = 8191s ;
  		etp_mf_fold_mir_bkhd_ct:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string etp_mf_fold_mir_bkhd_ct:coordinates = "start_of_scan_time" ;
  		string etp_mf_fold_mir_bkhd_ct:long_name = "Fold Mirror Bulkhead Center Temperature (Thermistor 6)" ;
  		string etp_mf_fold_mir_bkhd_ct:source = "APID826:ETP_MF_FOLD_MIR_BKHD_CT" ;
  	short etp_mf_ham_blkhd(scans) ;
  		etp_mf_ham_blkhd:_FillValue = -998s ;
  		etp_mf_ham_blkhd:valid_min = -8192s ;
  		etp_mf_ham_blkhd:valid_max = 8191s ;
  		etp_mf_ham_blkhd:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string etp_mf_ham_blkhd:coordinates = "start_of_scan_time" ;
  		string etp_mf_ham_blkhd:long_name = "Half-Angle Mirror Bulkhead Temperature (Thermistor 43)" ;
  		string etp_mf_ham_blkhd:source = "APID826:ETP_MF_HAM_BLKHD" ;
  	short etp_mf_km1_nxny(scans) ;
  		etp_mf_km1_nxny:_FillValue = -998s ;
  		etp_mf_km1_nxny:valid_min = -8192s ;
  		etp_mf_km1_nxny:valid_max = 8191s ;
  		etp_mf_km1_nxny:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string etp_mf_km1_nxny:coordinates = "start_of_scan_time" ;
  		string etp_mf_km1_nxny:long_name = "Kinematic Mount NX-NY Temperature (Thermistor 35)" ;
  		string etp_mf_km1_nxny:source = "APID826:ETP_MF_KM1_NXNY" ;
  	short etp_mf_km2_nxpy(scans) ;
  		etp_mf_km2_nxpy:_FillValue = -998s ;
  		etp_mf_km2_nxpy:valid_min = -8192s ;
  		etp_mf_km2_nxpy:valid_max = 8191s ;
  		etp_mf_km2_nxpy:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string etp_mf_km2_nxpy:coordinates = "start_of_scan_time" ;
  		string etp_mf_km2_nxpy:long_name = "Kinematic Mount NX-PY Temperature (Thermistor 34)" ;
  		string etp_mf_km2_nxpy:source = "APID826:ETP_MF_KM2_NXPY" ;
  	short etp_mf_km1_pxny(scans) ;
  		etp_mf_km1_pxny:_FillValue = -998s ;
  		etp_mf_km1_pxny:valid_min = -8192s ;
  		etp_mf_km1_pxny:valid_max = 8191s ;
  		etp_mf_km1_pxny:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string etp_mf_km1_pxny:coordinates = "start_of_scan_time" ;
  		string etp_mf_km1_pxny:long_name = "Kinematic Mount PX-NY Temperature (Thermistor 36)" ;
  		string etp_mf_km1_pxny:source = "APID826:ETP_MF_KM1_PXNY" ;
  	short etp_mf_km2_pxpy(scans) ;
  		etp_mf_km2_pxpy:_FillValue = -998s ;
  		etp_mf_km2_pxpy:valid_min = -8192s ;
  		etp_mf_km2_pxpy:valid_max = 8191s ;
  		etp_mf_km2_pxpy:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string etp_mf_km2_pxpy:coordinates = "start_of_scan_time" ;
  		string etp_mf_km2_pxpy:long_name = "Kinematic Mount PX-PY Temperature (Thermistor 37)" ;
  		string etp_mf_km2_pxpy:source = "APID826:ETP_MF_KM2_PXPY" ;
  	short etp_mf_nadir_raditr_nxp(scans) ;
  		etp_mf_nadir_raditr_nxp:_FillValue = -998s ;
  		etp_mf_nadir_raditr_nxp:valid_min = -8192s ;
  		etp_mf_nadir_raditr_nxp:valid_max = 8191s ;
  		etp_mf_nadir_raditr_nxp:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string etp_mf_nadir_raditr_nxp:coordinates = "start_of_scan_time" ;
  		string etp_mf_nadir_raditr_nxp:long_name = "Nadir Radiator NX-PY Temperature (Thermistor 15)" ;
  		string etp_mf_nadir_raditr_nxp:source = "APID826:ETP_MF_NADIR_RADITR_NXP" ;
  	short etp_mf_nadir_raditr_pxn(scans) ;
  		etp_mf_nadir_raditr_pxn:_FillValue = -998s ;
  		etp_mf_nadir_raditr_pxn:valid_min = -8192s ;
  		etp_mf_nadir_raditr_pxn:valid_max = 8191s ;
  		etp_mf_nadir_raditr_pxn:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string etp_mf_nadir_raditr_pxn:coordinates = "start_of_scan_time" ;
  		string etp_mf_nadir_raditr_pxn:long_name = "Nadir Radiator PX-NY Temperature (Thermistor 5)" ;
  		string etp_mf_nadir_raditr_pxn:source = "APID826:ETP_MF_NADIR_RADITR_PXN" ;
  	short etp_mf_scan_cavity_nx_n(scans) ;
  		etp_mf_scan_cavity_nx_n:_FillValue = -998s ;
  		etp_mf_scan_cavity_nx_n:valid_min = -8192s ;
  		etp_mf_scan_cavity_nx_n:valid_max = 8191s ;
  		etp_mf_scan_cavity_nx_n:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string etp_mf_scan_cavity_nx_n:coordinates = "start_of_scan_time" ;
  		string etp_mf_scan_cavity_nx_n:long_name = "Scan Cavity NX-NZ Temperature (Thermistor 47)" ;
  		string etp_mf_scan_cavity_nx_n:source = "APID826:ETP_MF_SCAN_CAVITY_NX_N" ;
  	short etp_mf_scan_cavity_nx_p(scans) ;
  		etp_mf_scan_cavity_nx_p:_FillValue = -998s ;
  		etp_mf_scan_cavity_nx_p:valid_min = -8192s ;
  		etp_mf_scan_cavity_nx_p:valid_max = 8191s ;
  		etp_mf_scan_cavity_nx_p:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string etp_mf_scan_cavity_nx_p:coordinates = "start_of_scan_time" ;
  		string etp_mf_scan_cavity_nx_p:long_name = "Scan Cavity NX-PZ Temperature (Thermistor 46)" ;
  		string etp_mf_scan_cavity_nx_p:source = "APID826:ETP_MF_SCAN_CAVITY_NX_P" ;
  	short etp_mf_scan_cvty_baf_nz(scans) ;
  		etp_mf_scan_cvty_baf_nz:_FillValue = -998s ;
  		etp_mf_scan_cvty_baf_nz:valid_min = -8192s ;
  		etp_mf_scan_cvty_baf_nz:valid_max = 8191s ;
  		etp_mf_scan_cvty_baf_nz:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string etp_mf_scan_cvty_baf_nz:coordinates = "start_of_scan_time" ;
  		string etp_mf_scan_cvty_baf_nz:long_name = "Scan Cavity Baffle NZ Temperature (Thermistor 10)" ;
  		string etp_mf_scan_cvty_baf_nz:source = "APID826:ETP_MF_SCAN_CVTY_BAF_NZ" ;
  	short etp_mf_scan_cvty_baf_pz(scans) ;
  		etp_mf_scan_cvty_baf_pz:_FillValue = -998s ;
  		etp_mf_scan_cvty_baf_pz:valid_min = -8192s ;
  		etp_mf_scan_cvty_baf_pz:valid_max = 8191s ;
  		etp_mf_scan_cvty_baf_pz:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string etp_mf_scan_cvty_baf_pz:coordinates = "start_of_scan_time" ;
  		string etp_mf_scan_cvty_baf_pz:long_name = "Scan Cavity Baffle PZ Temperature (Thermistor 9)" ;
  		string etp_mf_scan_cvty_baf_pz:source = "APID826:ETP_MF_SCAN_CVTY_BAF_PZ" ;
  	short etp_mf_scan_cvty_bkhd_n(scans) ;
  		etp_mf_scan_cvty_bkhd_n:_FillValue = -998s ;
  		etp_mf_scan_cvty_bkhd_n:valid_min = -8192s ;
  		etp_mf_scan_cvty_bkhd_n:valid_max = 8191s ;
  		etp_mf_scan_cvty_bkhd_n:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string etp_mf_scan_cvty_bkhd_n:coordinates = "start_of_scan_time" ;
  		string etp_mf_scan_cvty_bkhd_n:long_name = "Scan Cavity Bulkhead NY Temperature (Thermistor 8)" ;
  		string etp_mf_scan_cvty_bkhd_n:source = "APID826:ETP_MF_SCAN_CVTY_BKHD_N" ;
  	short etp_mf_space_radiator_n(scans) ;
  		etp_mf_space_radiator_n:_FillValue = -998s ;
  		etp_mf_space_radiator_n:valid_min = -8192s ;
  		etp_mf_space_radiator_n:valid_max = 8191s ;
  		etp_mf_space_radiator_n:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string etp_mf_space_radiator_n:coordinates = "start_of_scan_time" ;
  		string etp_mf_space_radiator_n:long_name = "Space Radiator NZ Temperature (Thermistor 41)" ;
  		string etp_mf_space_radiator_n:source = "APID826:ETP_MF_SPACE_RADIATOR_N" ;
  	short etp_mf_space_radiator_p(scans) ;
  		etp_mf_space_radiator_p:_FillValue = -998s ;
  		etp_mf_space_radiator_p:valid_min = -8192s ;
  		etp_mf_space_radiator_p:valid_max = 8191s ;
  		etp_mf_space_radiator_p:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string etp_mf_space_radiator_p:coordinates = "start_of_scan_time" ;
  		string etp_mf_space_radiator_p:long_name = "Space Radiator PZ Temperature (Thermistor 42)" ;
  		string etp_mf_space_radiator_p:source = "APID826:ETP_MF_SPACE_RADIATOR_P" ;
  	short etp_mf_stopassy_baff_nz(scans) ;
  		etp_mf_stopassy_baff_nz:_FillValue = -998s ;
  		etp_mf_stopassy_baff_nz:valid_min = -8192s ;
  		etp_mf_stopassy_baff_nz:valid_max = 8191s ;
  		etp_mf_stopassy_baff_nz:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string etp_mf_stopassy_baff_nz:coordinates = "start_of_scan_time" ;
  		string etp_mf_stopassy_baff_nz:long_name = "Aperture Stop Assembly Baffle NZ Temperature (Thermistor 14)" ;
  		string etp_mf_stopassy_baff_nz:source = "APID826:ETP_MF_STOPASSY_BAFF_NZ" ;
  	short etp_mf_tel_blkhd_nypz(scans) ;
  		etp_mf_tel_blkhd_nypz:_FillValue = -998s ;
  		etp_mf_tel_blkhd_nypz:valid_min = -8192s ;
  		etp_mf_tel_blkhd_nypz:valid_max = 8191s ;
  		etp_mf_tel_blkhd_nypz:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string etp_mf_tel_blkhd_nypz:coordinates = "start_of_scan_time" ;
  		string etp_mf_tel_blkhd_nypz:long_name = "Telescope Bulkhead NY-PZ Temperature (Thermistor 11)" ;
  		string etp_mf_tel_blkhd_nypz:source = "APID826:ETP_MF_TEL_BLKHD_NYPZ" ;
  	short etp_mf_tel_blkhd_py(scans) ;
  		etp_mf_tel_blkhd_py:_FillValue = -998s ;
  		etp_mf_tel_blkhd_py:valid_min = -8192s ;
  		etp_mf_tel_blkhd_py:valid_max = 8191s ;
  		etp_mf_tel_blkhd_py:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string etp_mf_tel_blkhd_py:coordinates = "start_of_scan_time" ;
  		string etp_mf_tel_blkhd_py:long_name = "Telescope Bulkhead PY Temperature (Thermistor 33)" ;
  		string etp_mf_tel_blkhd_py:source = "APID826:ETP_MF_TEL_BLKHD_PY" ;
  	short etp_se_a_hammtr_dfbear(scans) ;
  		etp_se_a_hammtr_dfbear:_FillValue = -998s ;
  		etp_se_a_hammtr_dfbear:valid_min = -8192s ;
  		etp_se_a_hammtr_dfbear:valid_max = 8191s ;
  		etp_se_a_hammtr_dfbear:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string etp_se_a_hammtr_dfbear:coordinates = "start_of_scan_time" ;
  		string etp_se_a_hammtr_dfbear:long_name = "SCE-A Half-Angle Mirror DF Bearing Motor Temperature (Thermistor 29)" ;
  		string etp_se_a_hammtr_dfbear:source = "APID826:ETP_SE_A_HAMMTR_DFBEAR" ;
  	short etp_se_a_telemtr_dfbear(scans) ;
  		etp_se_a_telemtr_dfbear:_FillValue = -998s ;
  		etp_se_a_telemtr_dfbear:valid_min = -8192s ;
  		etp_se_a_telemtr_dfbear:valid_max = 8191s ;
  		etp_se_a_telemtr_dfbear:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string etp_se_a_telemtr_dfbear:coordinates = "start_of_scan_time" ;
  		string etp_se_a_telemtr_dfbear:long_name = "SCE-A Telescope DF Bearing Motor Temperature (Thermistor 28)" ;
  		string etp_se_a_telemtr_dfbear:source = "APID826:ETP_SE_A_TELEMTR_DFBEAR" ;
  	short etp_se_b_hammtr_dfbear(scans) ;
  		etp_se_b_hammtr_dfbear:_FillValue = -998s ;
  		etp_se_b_hammtr_dfbear:valid_min = -8192s ;
  		etp_se_b_hammtr_dfbear:valid_max = 8191s ;
  		etp_se_b_hammtr_dfbear:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string etp_se_b_hammtr_dfbear:coordinates = "start_of_scan_time" ;
  		string etp_se_b_hammtr_dfbear:long_name = "SCE-B Half-Angle Mirror DF Bearing Motor Temperature (Thermistor 10)" ;
  		string etp_se_b_hammtr_dfbear:source = "APID826:ETP_SE_B_HAMMTR_DFBEAR" ;
  	short etp_se_b_telemtr_dfbear(scans) ;
  		etp_se_b_telemtr_dfbear:_FillValue = -998s ;
  		etp_se_b_telemtr_dfbear:valid_min = -8192s ;
  		etp_se_b_telemtr_dfbear:valid_max = 8191s ;
  		etp_se_b_telemtr_dfbear:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string etp_se_b_telemtr_dfbear:coordinates = "start_of_scan_time" ;
  		string etp_se_b_telemtr_dfbear:long_name = "SCE-B Telescope DF Bearing Motor Temperature (Thermistor 9)" ;
  		string etp_se_b_telemtr_dfbear:source = "APID826:ETP_SE_B_TELEMTR_DFBEAR" ;
  	short etp_ap_lw_cca(scans) ;
  		etp_ap_lw_cca:_FillValue = -998s ;
  		etp_ap_lw_cca:valid_min = -8192s ;
  		etp_ap_lw_cca:valid_max = 8191s ;
  		etp_ap_lw_cca:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string etp_ap_lw_cca:coordinates = "start_of_scan_time" ;
  		string etp_ap_lw_cca:long_name = "LW-IR Primary Circuit Card Assembly Temperature (Thermistor 1)" ;
  		string etp_ap_lw_cca:source = "APID826:ETP_AP_LW_CCA" ;
  	short etp_ap_sm_cca(scans) ;
  		etp_ap_sm_cca:_FillValue = -998s ;
  		etp_ap_sm_cca:valid_min = -8192s ;
  		etp_ap_sm_cca:valid_max = 8191s ;
  		etp_ap_sm_cca:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string etp_ap_sm_cca:coordinates = "start_of_scan_time" ;
  		string etp_ap_sm_cca:long_name = "SW/MW-IR Circuit Card Assembly Temperature (Thermistor 2)" ;
  		string etp_ap_sm_cca:source = "APID826:ETP_AP_SM_CCA" ;
  	short etp_ap_vn_cca(scans) ;
  		etp_ap_vn_cca:_FillValue = -998s ;
  		etp_ap_vn_cca:valid_min = -8192s ;
  		etp_ap_vn_cca:valid_max = 8191s ;
  		etp_ap_vn_cca:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string etp_ap_vn_cca:coordinates = "start_of_scan_time" ;
  		string etp_ap_vn_cca:long_name = "Visible/NIR Circuit Card Assembly Temperature (Thermistor 3)" ;
  		string etp_ap_vn_cca:source = "APID826:ETP_AP_VN_CCA" ;
  	short etp_dp_dnb_cca(scans) ;
  		etp_dp_dnb_cca:_FillValue = -998s ;
  		etp_dp_dnb_cca:valid_min = -8192s ;
  		etp_dp_dnb_cca:valid_max = 8191s ;
  		etp_dp_dnb_cca:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string etp_dp_dnb_cca:coordinates = "start_of_scan_time" ;
  		string etp_dp_dnb_cca:long_name = "Day/Night Band Circuit Card Assembly Temperature (Thermistor 60)" ;
  		string etp_dp_dnb_cca:source = "APID826:ETP_DP_DNB_CCA" ;
  	short etp_dp_dpp_cca(scans) ;
  		etp_dp_dpp_cca:_FillValue = -998s ;
  		etp_dp_dpp_cca:valid_min = -8192s ;
  		etp_dp_dpp_cca:valid_max = 8191s ;
  		etp_dp_dpp_cca:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string etp_dp_dpp_cca:coordinates = "start_of_scan_time" ;
  		string etp_dp_dpp_cca:long_name = "Digital Preprocessor Circuit Card Assembly Temperature (Thermistor 61)" ;
  		string etp_dp_dpp_cca:source = "APID826:ETP_DP_DPP_CCA" ;
  	short etp_dp_fpie_ad_cca(scans) ;
  		etp_dp_fpie_ad_cca:_FillValue = -998s ;
  		etp_dp_fpie_ad_cca:valid_min = -8192s ;
  		etp_dp_fpie_ad_cca:valid_max = 8191s ;
  		etp_dp_fpie_ad_cca:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string etp_dp_fpie_ad_cca:coordinates = "start_of_scan_time" ;
  		string etp_dp_fpie_ad_cca:long_name = "Focal Plane Integrated Electronics A/D Circuit Card Assembly Temperature (Thermistor 13)" ;
  		string etp_dp_fpie_ad_cca:source = "APID826:ETP_DP_FPIE_AD_CCA" ;
  	short etp_dp_fpie_clk_cca(scans) ;
  		etp_dp_fpie_clk_cca:_FillValue = -998s ;
  		etp_dp_fpie_clk_cca:valid_min = -8192s ;
  		etp_dp_fpie_clk_cca:valid_max = 8191s ;
  		etp_dp_fpie_clk_cca:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string etp_dp_fpie_clk_cca:coordinates = "start_of_scan_time" ;
  		string etp_dp_fpie_clk_cca:long_name = "Focal Plane Integrated Electronics Clock Circuit Card Assembly Temperature (Thermistor 51)" ;
  		string etp_dp_fpie_clk_cca:source = "APID826:ETP_DP_FPIE_CLK_CCA" ;
  	short etp_ft_cca(scans) ;
  		etp_ft_cca:_FillValue = -998s ;
  		etp_ft_cca:valid_min = -8192s ;
  		etp_ft_cca:valid_max = 8191s ;
  		etp_ft_cca:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string etp_ft_cca:coordinates = "start_of_scan_time" ;
  		string etp_ft_cca:long_name = "Focal Plane Temperature Controller Circuit Card Assembly Temperature (Thermistor 7)" ;
  		string etp_ft_cca:source = "APID826:ETP_FT_CCA" ;
  	short etp_ps1(scans) ;
  		etp_ps1:_FillValue = -998s ;
  		etp_ps1:valid_min = -8192s ;
  		etp_ps1:valid_max = 8191s ;
  		etp_ps1:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string etp_ps1:coordinates = "start_of_scan_time" ;
  		string etp_ps1:long_name = "Power Supply 1 Temperature (Thermistor 52)" ;
  		string etp_ps1:source = "APID826:ETP_PS1" ;
  	short etp_ps2(scans) ;
  		etp_ps2:_FillValue = -998s ;
  		etp_ps2:valid_min = -8192s ;
  		etp_ps2:valid_max = 8191s ;
  		etp_ps2:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string etp_ps2:coordinates = "start_of_scan_time" ;
  		string etp_ps2:long_name = "Power Supply 2 Temperature (Thermistor 53)" ;
  		string etp_ps2:source = "APID826:ETP_PS2" ;
  	short etp_se_a_cca(scans) ;
  		etp_se_a_cca:_FillValue = -998s ;
  		etp_se_a_cca:valid_min = -8192s ;
  		etp_se_a_cca:valid_max = 8191s ;
  		etp_se_a_cca:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string etp_se_a_cca:coordinates = "start_of_scan_time" ;
  		string etp_se_a_cca:long_name = "SCE-A Circuit Card Assembly Temperature (Thermistor 31)" ;
  		string etp_se_a_cca:source = "APID826:ETP_SE_A_CCA" ;
  	short etp_se_b_cca(scans) ;
  		etp_se_b_cca:_FillValue = -998s ;
  		etp_se_b_cca:valid_min = -8192s ;
  		etp_se_b_cca:valid_max = 8191s ;
  		etp_se_b_cca:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string etp_se_b_cca:coordinates = "start_of_scan_time" ;
  		string etp_se_b_cca:long_name = "SCE-B Circuit Card Assembly Temperature (Thermistor 12)" ;
  		string etp_se_b_cca:source = "APID826:ETP_SE_B_CCA" ;
  	ubyte ec_ft_lw_80k_setpt(scans) ;
  		ec_ft_lw_80k_setpt:_FillValue = 254UB ;
  		ec_ft_lw_80k_setpt:valid_min = 0UB ;
  		ec_ft_lw_80k_setpt:valid_max = 1UB ;
  		ec_ft_lw_80k_setpt:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string ec_ft_lw_80k_setpt:coordinates = "start_of_scan_time" ;
  		string ec_ft_lw_80k_setpt:long_name = "LW-IR 80K Setpoint Status" ;
  		string ec_ft_lw_80k_setpt:source = "APID826:EC_FT_LW_80K_SETPT" ;
  	ubyte ec_ft_lw_82k_setpt(scans) ;
  		ec_ft_lw_82k_setpt:_FillValue = 254UB ;
  		ec_ft_lw_82k_setpt:valid_min = 0UB ;
  		ec_ft_lw_82k_setpt:valid_max = 1UB ;
  		ec_ft_lw_82k_setpt:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string ec_ft_lw_82k_setpt:coordinates = "start_of_scan_time" ;
  		string ec_ft_lw_82k_setpt:long_name = "LW-IR 82K Setpoint Status" ;
  		string ec_ft_lw_82k_setpt:source = "APID826:EC_FT_LW_82K_SETPT" ;
  	ubyte ec_ft_sm_80k_setpt(scans) ;
  		ec_ft_sm_80k_setpt:_FillValue = 254UB ;
  		ec_ft_sm_80k_setpt:valid_min = 0UB ;
  		ec_ft_sm_80k_setpt:valid_max = 1UB ;
  		ec_ft_sm_80k_setpt:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string ec_ft_sm_80k_setpt:coordinates = "start_of_scan_time" ;
  		string ec_ft_sm_80k_setpt:long_name = "SW/MW-IR 80K Setpoint Status" ;
  		string ec_ft_sm_80k_setpt:source = "APID826:EC_FT_SM_80K_SETPT" ;
  	ubyte ec_ft_sm_82k_setpt(scans) ;
  		ec_ft_sm_82k_setpt:_FillValue = 254UB ;
  		ec_ft_sm_82k_setpt:valid_min = 0UB ;
  		ec_ft_sm_82k_setpt:valid_max = 1UB ;
  		ec_ft_sm_82k_setpt:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string ec_ft_sm_82k_setpt:coordinates = "start_of_scan_time" ;
  		string ec_ft_sm_82k_setpt:long_name = "SW/MW-IR 82K Setpoint Status" ;
  		string ec_ft_sm_82k_setpt:source = "APID826:EC_FT_SM_82K_SETPT" ;
  	ubyte ec_ft_lw_htr_on(scans) ;
  		ec_ft_lw_htr_on:_FillValue = 254UB ;
  		ec_ft_lw_htr_on:valid_min = 0UB ;
  		ec_ft_lw_htr_on:valid_max = 1UB ;
  		ec_ft_lw_htr_on:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string ec_ft_lw_htr_on:coordinates = "start_of_scan_time" ;
  		string ec_ft_lw_htr_on:long_name = "LW-IR Heater Status" ;
  		string ec_ft_lw_htr_on:source = "APID826:EC_FT_LW_HTR_ON" ;
  	ubyte ec_ft_sm_htr_on(scans) ;
  		ec_ft_sm_htr_on:_FillValue = 254UB ;
  		ec_ft_sm_htr_on:valid_min = 0UB ;
  		ec_ft_sm_htr_on:valid_max = 1UB ;
  		ec_ft_sm_htr_on:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string ec_ft_sm_htr_on:coordinates = "start_of_scan_time" ;
  		string ec_ft_sm_htr_on:long_name = "SW/MW-IR Heater Status" ;
  		string ec_ft_sm_htr_on:source = "APID826:EC_FT_SM_HTR_ON" ;
  	ubyte ec_hm_dnb_htr_cntl(scans) ;
  		ec_hm_dnb_htr_cntl:_FillValue = 254UB ;
  		ec_hm_dnb_htr_cntl:valid_min = 0UB ;
  		ec_hm_dnb_htr_cntl:valid_max = 1UB ;
  		ec_hm_dnb_htr_cntl:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string ec_hm_dnb_htr_cntl:coordinates = "start_of_scan_time" ;
  		string ec_hm_dnb_htr_cntl:long_name = "Day/Night Band Heater Control Echo" ;
  		string ec_hm_dnb_htr_cntl:source = "APID826:EC_HM_DNB_HTR_CNTL" ;
  	ubyte ec_hm_ham_op_htr_cntl(scans) ;
  		ec_hm_ham_op_htr_cntl:_FillValue = 254UB ;
  		ec_hm_ham_op_htr_cntl:valid_min = 0UB ;
  		ec_hm_ham_op_htr_cntl:valid_max = 1UB ;
  		ec_hm_ham_op_htr_cntl:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string ec_hm_ham_op_htr_cntl:coordinates = "start_of_scan_time" ;
  		string ec_hm_ham_op_htr_cntl:long_name = "Half-Angle Mirror Control Echo" ;
  		string ec_hm_ham_op_htr_cntl:source = "APID826:EC_HM_HAM_OP_HTR_CNTL" ;
  	ubyte ec_hm_tel_op_htr_cntl(scans) ;
  		ec_hm_tel_op_htr_cntl:_FillValue = 254UB ;
  		ec_hm_tel_op_htr_cntl:valid_min = 0UB ;
  		ec_hm_tel_op_htr_cntl:valid_max = 1UB ;
  		ec_hm_tel_op_htr_cntl:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string ec_hm_tel_op_htr_cntl:coordinates = "start_of_scan_time" ;
  		string ec_hm_tel_op_htr_cntl:long_name = "Telescope Operational Heater Control Echo" ;
  		string ec_hm_tel_op_htr_cntl:source = "APID826:EC_HM_TEL_OP_HTR_CNTL" ;
  	ushort ec_hm_ham_ophtr_temp_se(scans) ;
  		ec_hm_ham_ophtr_temp_se:_FillValue = 65534US ;
  		ec_hm_ham_ophtr_temp_se:valid_min = 0US ;
  		ec_hm_ham_ophtr_temp_se:valid_max = 16383US ;
  		ec_hm_ham_ophtr_temp_se:missing_value = 65528US, 65529US, 65530US, 65531US, 65532US, 65533US, 65534US, 65535US ;
  		string ec_hm_ham_ophtr_temp_se:coordinates = "start_of_scan_time" ;
  		string ec_hm_ham_ophtr_temp_se:long_name = "Half-Angle Mirror Operational Heater Setpoint Echo" ;
  		string ec_hm_ham_ophtr_temp_se:source = "APID826:EC_HM_HAM_OPHTR_TEMP_SE" ;
  	ushort ec_hm_tel_ophtr_temp_set(scans) ;
  		ec_hm_tel_ophtr_temp_set:_FillValue = 65534US ;
  		ec_hm_tel_ophtr_temp_set:valid_min = 0US ;
  		ec_hm_tel_ophtr_temp_set:valid_max = 16383US ;
  		ec_hm_tel_ophtr_temp_set:missing_value = 65528US, 65529US, 65530US, 65531US, 65532US, 65533US, 65534US, 65535US ;
  		string ec_hm_tel_ophtr_temp_set:coordinates = "start_of_scan_time" ;
  		string ec_hm_tel_ophtr_temp_set:long_name = "Telescope Operational Heater Setpoint Echo" ;
  		string ec_hm_tel_ophtr_temp_set:source = "APID826:EC_HM_TEL_OPHTR_TEMP_SET" ;
  	ushort etp_bb_avg_temp(scans) ;
  		etp_bb_avg_temp:_FillValue = 65534US ;
  		etp_bb_avg_temp:valid_min = 0US ;
  		etp_bb_avg_temp:valid_max = 16383US ;
  		etp_bb_avg_temp:missing_value = 65528US, 65529US, 65530US, 65531US, 65532US, 65533US, 65534US, 65535US ;
  		string etp_bb_avg_temp:coordinates = "start_of_scan_time" ;
  		string etp_bb_avg_temp:long_name = "Blackbody Average Temperature" ;
  		string etp_bb_avg_temp:source = "APID826:ETP_BB_AVG_TEMP" ;
  	ushort ec_bb_htr_temp_set(scans) ;
  		ec_bb_htr_temp_set:_FillValue = 65534US ;
  		ec_bb_htr_temp_set:valid_min = 0US ;
  		ec_bb_htr_temp_set:valid_max = 16383US ;
  		ec_bb_htr_temp_set:missing_value = 65528US, 65529US, 65530US, 65531US, 65532US, 65533US, 65534US, 65535US ;
  		string ec_bb_htr_temp_set:coordinates = "start_of_scan_time" ;
  		string ec_bb_htr_temp_set:long_name = "Blackbody Heater Temperature Setpoint Echo" ;
  		string ec_bb_htr_temp_set:source = "APID826:EC_BB_HTR_TEMP_SET" ;
  	ushort ec_bb_select(scans) ;
  		ec_bb_select:_FillValue = 65534US ;
  		ec_bb_select:valid_min = 0US ;
  		ec_bb_select:valid_max = 65535US ;
  		ec_bb_select:missing_value = 65528US, 65529US, 65530US, 65531US, 65532US, 65533US, 65534US, 65535US ;
  		string ec_bb_select:coordinates = "start_of_scan_time" ;
  		string ec_bb_select:long_name = "Blackbody Average Temperature Thermistor Select Status" ;
  		string ec_bb_select:source = "APID826:EC_BB_SELECT" ;
  	ubyte s_sd_position(scans) ;
  		s_sd_position:_FillValue = 254UB ;
  		s_sd_position:valid_min = 0UB ;
  		s_sd_position:valid_max = 255UB ;
  		s_sd_position:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string s_sd_position:coordinates = "start_of_scan_time" ;
  		string s_sd_position:long_name = "SDSM  Position" ;
  		string s_sd_position:source = "APID826:S_SD_POSITION" ;
  	short v_sd_sdsm_amp_samples(scans, sdsm_detectors_750m, sdsm_samples) ;
  		v_sd_sdsm_amp_samples:_FillValue = -998s ;
  		v_sd_sdsm_amp_samples:valid_min = -8192s ;
  		v_sd_sdsm_amp_samples:valid_max = 8191s ;
  		v_sd_sdsm_amp_samples:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string v_sd_sdsm_amp_samples:coordinates = "start_of_scan_time" ;
  		string v_sd_sdsm_amp_samples:long_name = "SDSM  Amp Sample Voltages" ;
  		string v_sd_sdsm_amp_samples:source = "APID826:V_SD_SDSM_AMP1-8_SMPL1-5" ;
  	short etp_sd_sdsm_preamp(scans) ;
  		etp_sd_sdsm_preamp:_FillValue = -998s ;
  		etp_sd_sdsm_preamp:valid_min = -8192s ;
  		etp_sd_sdsm_preamp:valid_max = 8191s ;
  		etp_sd_sdsm_preamp:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string etp_sd_sdsm_preamp:coordinates = "start_of_scan_time" ;
  		string etp_sd_sdsm_preamp:long_name = "SDSM PreAmp Temperature (Thermistor 57)" ;
  		string etp_sd_sdsm_preamp:source = "APID826:ETP_SD_SDSM_PREAMP" ;
  	ubyte ec_sd_sdsm_mtr_hold(scans) ;
  		ec_sd_sdsm_mtr_hold:_FillValue = 254UB ;
  		ec_sd_sdsm_mtr_hold:valid_min = 0UB ;
  		ec_sd_sdsm_mtr_hold:valid_max = 1UB ;
  		ec_sd_sdsm_mtr_hold:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string ec_sd_sdsm_mtr_hold:coordinates = "start_of_scan_time" ;
  		string ec_sd_sdsm_mtr_hold:long_name = "SDSM Motor Hold Status" ;
  		string ec_sd_sdsm_mtr_hold:source = "APID826:EC_SD_SDSM_MTR_HOLD" ;
  	ubyte ec_sd_preamp_even_pwr(scans) ;
  		ec_sd_preamp_even_pwr:_FillValue = 254UB ;
  		ec_sd_preamp_even_pwr:valid_min = 0UB ;
  		ec_sd_preamp_even_pwr:valid_max = 1UB ;
  		ec_sd_preamp_even_pwr:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string ec_sd_preamp_even_pwr:coordinates = "start_of_scan_time" ;
  		string ec_sd_preamp_even_pwr:long_name = "SDSM PreAmp 2,4,6,8 Power Status" ;
  		string ec_sd_preamp_even_pwr:source = "APID826:EC_SD_PREAMP_EVEN_PWR" ;
  	ubyte ec_sd_preamp_odd_pwr(scans) ;
  		ec_sd_preamp_odd_pwr:_FillValue = 254UB ;
  		ec_sd_preamp_odd_pwr:valid_min = 0UB ;
  		ec_sd_preamp_odd_pwr:valid_max = 1UB ;
  		ec_sd_preamp_odd_pwr:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string ec_sd_preamp_odd_pwr:coordinates = "start_of_scan_time" ;
  		string ec_sd_preamp_odd_pwr:long_name = "SDSM PreAmp 1,3,5,7 Power Status" ;
  		string ec_sd_preamp_odd_pwr:source = "APID826:EC_SD_PREAMP_ODD_PWR" ;
  	ubyte ec_sd_sdsm_mtr_at_home(scans) ;
  		ec_sd_sdsm_mtr_at_home:_FillValue = 254UB ;
  		ec_sd_sdsm_mtr_at_home:valid_min = 0UB ;
  		ec_sd_sdsm_mtr_at_home:valid_max = 1UB ;
  		ec_sd_sdsm_mtr_at_home:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string ec_sd_sdsm_mtr_at_home:coordinates = "start_of_scan_time" ;
  		string ec_sd_sdsm_mtr_at_home:long_name = "SDSM Motor At Home Status" ;
  		string ec_sd_sdsm_mtr_at_home:source = "APID826:EC_SD_SDSM_MTR_AT_HOME" ;
  	ushort s_se_tele_timestmps(scans, encoder_samples) ;
  		s_se_tele_timestmps:_FillValue = 65534US ;
  		s_se_tele_timestmps:valid_min = 0US ;
  		s_se_tele_timestmps:valid_max = 65535US ;
  		s_se_tele_timestmps:missing_value = 65528US, 65529US, 65530US, 65531US, 65532US, 65533US, 65534US, 65535US ;
  		string s_se_tele_timestmps:coordinates = "start_of_scan_time" ;
  		string s_se_tele_timestmps:long_name = "Telescope Pulse Arrival Timestamps" ;
  		string s_se_tele_timestmps:source = "APID826:S_SE_TELE_TIMESTMP_0000-1289" ;
  	ushort s_se_ham_timestmps(scans, encoder_samples) ;
  		s_se_ham_timestmps:_FillValue = 65534US ;
  		s_se_ham_timestmps:valid_min = 0US ;
  		s_se_ham_timestmps:valid_max = 65535US ;
  		s_se_ham_timestmps:missing_value = 65528US, 65529US, 65530US, 65531US, 65532US, 65533US, 65534US, 65535US ;
  		string s_se_ham_timestmps:coordinates = "start_of_scan_time" ;
  		string s_se_ham_timestmps:long_name = "Half-Angle Mirror Pulse Arrival Timestamps" ;
  		string s_se_ham_timestmps:source = "APID826:S_SE_HAM_TIMESTMP_0000-1289" ;
  	ushort s_dp_tele_ang_scan_strt(scans) ;
  		s_dp_tele_ang_scan_strt:_FillValue = 65534US ;
  		s_dp_tele_ang_scan_strt:valid_min = 0US ;
  		s_dp_tele_ang_scan_strt:valid_max = 65535US ;
  		s_dp_tele_ang_scan_strt:missing_value = 65528US, 65529US, 65530US, 65531US, 65532US, 65533US, 65534US, 65535US ;
  		string s_dp_tele_ang_scan_strt:coordinates = "start_of_scan_time" ;
  		string s_dp_tele_ang_scan_strt:long_name = "Telescope Raw Angle Count At Scan Start" ;
  		string s_dp_tele_ang_scan_strt:source = "APID826:S_DP_TELE_ANG_SCAN_STRT" ;
  	ushort s_dp_ham_ang_scan_strt(scans) ;
  		s_dp_ham_ang_scan_strt:_FillValue = 65534US ;
  		s_dp_ham_ang_scan_strt:valid_min = 0US ;
  		s_dp_ham_ang_scan_strt:valid_max = 65535US ;
  		s_dp_ham_ang_scan_strt:missing_value = 65528US, 65529US, 65530US, 65531US, 65532US, 65533US, 65534US, 65535US ;
  		string s_dp_ham_ang_scan_strt:coordinates = "start_of_scan_time" ;
  		string s_dp_ham_ang_scan_strt:long_name = "Half-Angle Mirror Raw Angle Count At Scan Start" ;
  		string s_dp_ham_ang_scan_strt:source = "APID826:S_DP_HAM_ANG_SCAN_STRT" ;
  	short es_cp_hrdt_values(scans, hrdt_samples) ;
  		es_cp_hrdt_values:_FillValue = -998s ;
  		es_cp_hrdt_values:valid_min = -8192s ;
  		es_cp_hrdt_values:valid_max = 8191s ;
  		es_cp_hrdt_values:missing_value = -992s, -993s, -994s, -995s, -996s, -997s, -998s, -999s ;
  		string es_cp_hrdt_values:coordinates = "start_of_scan_time" ;
  		string es_cp_hrdt_values:long_name = "Hi-Rate Dwell Telemetry Point Values" ;
  		string es_cp_hrdt_values:source = "APID826:ES_CP_HRDT_VALUE_1-16" ;
  	ushort c_cp_hrdt_muxaddr(scans) ;
  		c_cp_hrdt_muxaddr:_FillValue = 65534US ;
  		c_cp_hrdt_muxaddr:valid_min = 0US ;
  		c_cp_hrdt_muxaddr:valid_max = 65535US ;
  		c_cp_hrdt_muxaddr:missing_value = 65528US, 65529US, 65530US, 65531US, 65532US, 65533US, 65534US, 65535US ;
  		string c_cp_hrdt_muxaddr:coordinates = "start_of_scan_time" ;
  		string c_cp_hrdt_muxaddr:long_name = "Hi-Rate Dwell Telemetry Point Mux Address Selection" ;
  		string c_cp_hrdt_muxaddr:source = "APID826:C_CP_HRDT_MUXADDR" ;
  } // group Engineering_Data

group: Image_375m {
  dimensions:
  	band = 5 ;
  	line = UNLIMITED ; // (6144 currently)
  	pixel = 6400 ;
  	calib_source = 3 ;
  	cal_samples = 96 ;
  variables:
  	string band(band) ;
  		string band:long_name = "wavelength band identifier" ;
  	string calib_source(calib_source) ;
  		string calib_source:long_name = "calibration source identifier" ;
  	int lines_per_granule(granules) ;
  		lines_per_granule:_FillValue = -998 ;
  		lines_per_granule:valid_min = -2147483648 ;
  		lines_per_granule:valid_max = 2147483647 ;
  		lines_per_granule:missing_value = -992, -993, -994, -995, -996, -997, -998, -999 ;
  		string lines_per_granule:long_name = "Number of lines for each granule" ;
  	int starting_line_per_granule(granules) ;
  		starting_line_per_granule:_FillValue = -998 ;
  		starting_line_per_granule:valid_min = -2147483648 ;
  		starting_line_per_granule:valid_max = 2147483647 ;
  		starting_line_per_granule:missing_value = -992, -993, -994, -995, -996, -997, -998, -999 ;
  		string starting_line_per_granule:long_name = "Index of the line that starts each granule" ;
  	double earthview_start_of_data(band, scans) ;
  		earthview_start_of_data:_FillValue = -999.8 ;
  		earthview_start_of_data:valid_min = 1.48323e+15 ;
  		earthview_start_of_data:valid_max = 2.27215e+15 ;
  		earthview_start_of_data:missing_value = -999.2, -999.3, -999.4, -999.5, -999.6, -999.7, -999.8, -999.9 ;
  		string earthview_start_of_data:coordinates = "band" ;
  		string earthview_start_of_data:units = "microseconds since 1958/01/01 00:00:00" ;
  		string earthview_start_of_data:long_name = "Time at scan start" ;
  		string earthview_start_of_data:source = "(APID818, APID819, APID820, APID813, APID817):TimeOfDayStartOfData" ;
  		string earthview_start_of_data:standard_name = "time" ;
  	double earthview_scan_terminus(band, scans) ;
  		earthview_scan_terminus:_FillValue = -999.8 ;
  		earthview_scan_terminus:valid_min = 1.48323e+15 ;
  		earthview_scan_terminus:valid_max = 2.27215e+15 ;
  		earthview_scan_terminus:missing_value = -999.2, -999.3, -999.4, -999.5, -999.6, -999.7, -999.8, -999.9 ;
  		string earthview_scan_terminus:coordinates = "band" ;
  		string earthview_scan_terminus:units = "microseconds since 1958/01/01 00:00:00" ;
  		string earthview_scan_terminus:long_name = "Time at scan terminus" ;
  		string earthview_scan_terminus:source = "(APID818, APID819, APID820, APID813, APID817):ScanTerminus" ;
  		string earthview_scan_terminus:standard_name = "time" ;
  	double calibview_start_of_data(band, scans) ;
  		calibview_start_of_data:_FillValue = -999.8 ;
  		calibview_start_of_data:valid_min = 1.48323e+15 ;
  		calibview_start_of_data:valid_max = 2.27215e+15 ;
  		calibview_start_of_data:missing_value = -999.2, -999.3, -999.4, -999.5, -999.6, -999.7, -999.8, -999.9 ;
  		string calibview_start_of_data:coordinates = "band" ;
  		string calibview_start_of_data:units = "microseconds since 1958/01/01 00:00:00" ;
  		string calibview_start_of_data:long_name = "Time at scan start" ;
  		string calibview_start_of_data:source = "APID825:TimeOfDayStartOfData (for each included band)" ;
  		string calibview_start_of_data:standard_name = "time" ;
  	double calibview_scan_terminus(band, scans) ;
  		calibview_scan_terminus:_FillValue = -999.8 ;
  		calibview_scan_terminus:valid_min = 1.48323e+15 ;
  		calibview_scan_terminus:valid_max = 2.27215e+15 ;
  		calibview_scan_terminus:missing_value = -999.2, -999.3, -999.4, -999.5, -999.6, -999.7, -999.8, -999.9 ;
  		string calibview_scan_terminus:coordinates = "band" ;
  		string calibview_scan_terminus:units = "microseconds since 1958/01/01 00:00:00" ;
  		string calibview_scan_terminus:long_name = "Time at scan terminus" ;
  		string calibview_scan_terminus:source = "APID825:ScanTerminus (for each included band)" ;
  		string calibview_scan_terminus:standard_name = "time" ;
  	uint earthview_band_control_word(band, scans) ;
  		earthview_band_control_word:_FillValue = 4294967294U ;
  		earthview_band_control_word:valid_min = 0U ;
  		earthview_band_control_word:valid_max = 4294967295U ;
  		earthview_band_control_word:missing_value = 4294967288U, 0U, 4294967289U, 0U, 4294967290U, 0U, 4294967291U, 0U ;
  		string earthview_band_control_word:coordinates = "band earthview_start_of_data" ;
  		string earthview_band_control_word:long_name = "Earth view Band Control Word" ;
  		string earthview_band_control_word:source = "(APID818, APID819, APID820, APID813, APID817):BandControlWord" ;
  	uint calibview_band_control_word(band, scans) ;
  		calibview_band_control_word:_FillValue = 4294967294U ;
  		calibview_band_control_word:valid_min = 0U ;
  		calibview_band_control_word:valid_max = 4294967295U ;
  		calibview_band_control_word:missing_value = 4294967288U, 0U, 4294967289U, 0U, 4294967290U, 0U, 4294967291U, 0U ;
  		string calibview_band_control_word:coordinates = "band calibview_start_of_data" ;
  		string calibview_band_control_word:long_name = "Calibration view Band Control Word" ;
  		string calibview_band_control_word:source = "APID825:BandControlWord (for each included band)" ;
  	ushort earthview(band, line, pixel) ;
  		earthview:_FillValue = 65534US ;
  		earthview:valid_min = 0US ;
  		earthview:valid_max = 4095US ;
  		earthview:missing_value = 65528US, 65529US, 65530US, 65531US, 65532US, 65533US, 65534US, 65535US ;
  		string earthview:coordinates = "band earthview_start_of_data" ;
  		string earthview:long_name = "Digital counts from the Earth view for Image bands 1-5" ;
  		string earthview:source = "APID818, APID819, APID820, APID813, APID817" ;
  		earthview:chunk_size = 1, 6144, 6400 ;
  		earthview:chunk_compression_level = 2 ;
  	ushort calibview(band, calib_source, line, cal_samples) ;
  		calibview:_FillValue = 65534US ;
  		calibview:valid_min = 0US ;
  		calibview:valid_max = 16383US ;
  		calibview:missing_value = 65528US, 65529US, 65530US, 65531US, 65532US, 65533US, 65534US, 65535US ;
  		string calibview:coordinates = "band calib_source calibview_start_of_data" ;
  		string calibview:long_name = "Digital counts from the space view, black body, and solar diffuser for Image bands 1-5" ;
  		string calibview:source = "APID825" ;
  		calibview:chunk_size = 1, 3, 6144, 96 ;
  		calibview:chunk_compression_level = 2 ;
  } // group Image_375m

group: Image_750m_DualGain {
  dimensions:
  	band = 7 ;
  	line = UNLIMITED ; // (3072 currently)
  	pixel = 6304 ;
  	calib_source = 3 ;
  	cal_samples = 48 ;
  variables:
  	string band(band) ;
  		string band:long_name = "wavelength band identifier" ;
  	string calib_source(calib_source) ;
  		string calib_source:long_name = "calibration source identifier" ;
  	int lines_per_granule(granules) ;
  		lines_per_granule:_FillValue = -998 ;
  		lines_per_granule:valid_min = -2147483648 ;
  		lines_per_granule:valid_max = 2147483647 ;
  		lines_per_granule:missing_value = -992, -993, -994, -995, -996, -997, -998, -999 ;
  		string lines_per_granule:long_name = "Number of lines for each granule" ;
  	int starting_line_per_granule(granules) ;
  		starting_line_per_granule:_FillValue = -998 ;
  		starting_line_per_granule:valid_min = -2147483648 ;
  		starting_line_per_granule:valid_max = 2147483647 ;
  		starting_line_per_granule:missing_value = -992, -993, -994, -995, -996, -997, -998, -999 ;
  		string starting_line_per_granule:long_name = "Index of the line that starts each granule" ;
  	double earthview_start_of_data(band, scans) ;
  		earthview_start_of_data:_FillValue = -999.8 ;
  		earthview_start_of_data:valid_min = 1.48323e+15 ;
  		earthview_start_of_data:valid_max = 2.27215e+15 ;
  		earthview_start_of_data:missing_value = -999.2, -999.3, -999.4, -999.5, -999.6, -999.7, -999.8, -999.9 ;
  		string earthview_start_of_data:coordinates = "band" ;
  		string earthview_start_of_data:units = "microseconds since 1958/01/01 00:00:00" ;
  		string earthview_start_of_data:long_name = "Time at scan start" ;
  		string earthview_start_of_data:source = "(APID804, APID803, APID802, APID800, APID801, APID806, APID811):TimeOfDayStartOfData" ;
  		string earthview_start_of_data:standard_name = "time" ;
  	double earthview_scan_terminus(band, scans) ;
  		earthview_scan_terminus:_FillValue = -999.8 ;
  		earthview_scan_terminus:valid_min = 1.48323e+15 ;
  		earthview_scan_terminus:valid_max = 2.27215e+15 ;
  		earthview_scan_terminus:missing_value = -999.2, -999.3, -999.4, -999.5, -999.6, -999.7, -999.8, -999.9 ;
  		string earthview_scan_terminus:coordinates = "band" ;
  		string earthview_scan_terminus:units = "microseconds since 1958/01/01 00:00:00" ;
  		string earthview_scan_terminus:long_name = "Time at scan terminus" ;
  		string earthview_scan_terminus:source = "(APID804, APID803, APID802, APID800, APID801, APID806, APID811):ScanTerminus" ;
  		string earthview_scan_terminus:standard_name = "time" ;
  	double calibview_start_of_data(band, scans) ;
  		calibview_start_of_data:_FillValue = -999.8 ;
  		calibview_start_of_data:valid_min = 1.48323e+15 ;
  		calibview_start_of_data:valid_max = 2.27215e+15 ;
  		calibview_start_of_data:missing_value = -999.2, -999.3, -999.4, -999.5, -999.6, -999.7, -999.8, -999.9 ;
  		string calibview_start_of_data:coordinates = "band" ;
  		string calibview_start_of_data:units = "microseconds since 1958/01/01 00:00:00" ;
  		string calibview_start_of_data:long_name = "Time at scan start" ;
  		string calibview_start_of_data:source = "APID825:TimeOfDayStartOfData (for each included band)" ;
  		string calibview_start_of_data:standard_name = "time" ;
  	double calibview_scan_terminus(band, scans) ;
  		calibview_scan_terminus:_FillValue = -999.8 ;
  		calibview_scan_terminus:valid_min = 1.48323e+15 ;
  		calibview_scan_terminus:valid_max = 2.27215e+15 ;
  		calibview_scan_terminus:missing_value = -999.2, -999.3, -999.4, -999.5, -999.6, -999.7, -999.8, -999.9 ;
  		string calibview_scan_terminus:coordinates = "band" ;
  		string calibview_scan_terminus:units = "microseconds since 1958/01/01 00:00:00" ;
  		string calibview_scan_terminus:long_name = "Time at scan terminus" ;
  		string calibview_scan_terminus:source = "APID825:ScanTerminus (for each included band)" ;
  		string calibview_scan_terminus:standard_name = "time" ;
  	uint earthview_band_control_word(band, scans) ;
  		earthview_band_control_word:_FillValue = 4294967294U ;
  		earthview_band_control_word:valid_min = 0U ;
  		earthview_band_control_word:valid_max = 4294967295U ;
  		earthview_band_control_word:missing_value = 4294967288U, 0U, 4294967289U, 0U, 4294967290U, 0U, 4294967291U, 0U ;
  		string earthview_band_control_word:coordinates = "band earthview_start_of_data" ;
  		string earthview_band_control_word:long_name = "Earth view Band Control Word" ;
  		string earthview_band_control_word:source = "(APID804, APID803, APID802, APID800, APID801, APID806, APID811):BandControlWord" ;
  	uint calibview_band_control_word(band, scans) ;
  		calibview_band_control_word:_FillValue = 4294967294U ;
  		calibview_band_control_word:valid_min = 0U ;
  		calibview_band_control_word:valid_max = 4294967295U ;
  		calibview_band_control_word:missing_value = 4294967288U, 0U, 4294967289U, 0U, 4294967290U, 0U, 4294967291U, 0U ;
  		string calibview_band_control_word:coordinates = "band calibview_start_of_data" ;
  		string calibview_band_control_word:long_name = "Calibration view Band Control Word" ;
  		string calibview_band_control_word:source = "APID825:BandControlWord (for each included band)" ;
  	ushort earthview(band, line, pixel) ;
  		earthview:_FillValue = 65534US ;
  		earthview:valid_min = 0US ;
  		earthview:valid_max = 4095US ;
  		earthview:missing_value = 65528US, 65529US, 65530US, 65531US, 65532US, 65533US, 65534US, 65535US ;
  		string earthview:coordinates = "band earthview_start_of_data" ;
  		string earthview:long_name = "Digital counts from the Earth view for Moderate dual gain bands 1-5, 7, 13" ;
  		string earthview:source = "APID804, APID803, APID802, APID800, APID801, APID806, APID811" ;
  		earthview:chunk_size = 1, 3072, 6304 ;
  		earthview:chunk_compression_level = 2 ;
  	ubyte earthview_gain(band, line, pixel) ;
  		earthview_gain:_FillValue = 254UB ;
  		earthview_gain:valid_min = 0UB ;
  		earthview_gain:valid_max = 1UB ;
  		earthview_gain:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string earthview_gain:coordinates = "band earthview_start_of_data" ;
  		string earthview_gain:long_name = "Gain state from the Earth view for Moderate dual gain bands 1-5, 7, 13" ;
  		string earthview_gain:source = "APID804, APID803, APID802, APID800, APID801, APID806, APID811" ;
  		earthview_gain:chunk_size = 1, 3072, 6304 ;
  		earthview_gain:chunk_compression_level = 2 ;
  	ushort calibview(band, calib_source, line, cal_samples) ;
  		calibview:_FillValue = 65534US ;
  		calibview:valid_min = 0US ;
  		calibview:valid_max = 16383US ;
  		calibview:missing_value = 65528US, 65529US, 65530US, 65531US, 65532US, 65533US, 65534US, 65535US ;
  		string calibview:coordinates = "band calib_source calibview_start_of_data" ;
  		string calibview:long_name = "Digital counts from the space view, black body, and solar diffuser for Moderate dual gain bands 1-5, 7, 13" ;
  		string calibview:source = "APID825" ;
  		calibview:chunk_size = 1, 3, 3072, 48 ;
  		calibview:chunk_compression_level = 2 ;
  	ubyte calibview_gain(band, calib_source, line, cal_samples) ;
  		calibview_gain:_FillValue = 254UB ;
  		calibview_gain:valid_min = 0UB ;
  		calibview_gain:valid_max = 1UB ;
  		calibview_gain:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string calibview_gain:coordinates = "band calib_source calibview_start_of_data" ;
  		string calibview_gain:long_name = "Gain state from the space view, black body, and solar diffuser for Moderate dual gain bands 1-5, 7, 13" ;
  		string calibview_gain:source = "APID825" ;
  		calibview_gain:chunk_size = 1, 3, 3072, 48 ;
  		calibview_gain:chunk_compression_level = 2 ;
  } // group Image_750m_DualGain

group: Image_750m_SingleGain {
  dimensions:
  	band = 9 ;
  	line = UNLIMITED ; // (3072 currently)
  	pixel = 3200 ;
  	calib_band = 10 ;
  	calib_source = 3 ;
  	cal_samples = 48 ;
  variables:
  	string band(band) ;
  		string band:long_name = "earthview wavelength band identifier" ;
  	string calib_band(calib_band) ;
  		string calib_band:long_name = "calibration view wavelength band identifier" ;
  	string calib_source(calib_source) ;
  		string calib_source:long_name = "calibration source identifier" ;
  	int lines_per_granule(granules) ;
  		lines_per_granule:_FillValue = -998 ;
  		lines_per_granule:valid_min = -2147483648 ;
  		lines_per_granule:valid_max = 2147483647 ;
  		lines_per_granule:missing_value = -992, -993, -994, -995, -996, -997, -998, -999 ;
  		string lines_per_granule:long_name = "Number of lines for each granule" ;
  	int starting_line_per_granule(granules) ;
  		starting_line_per_granule:_FillValue = -998 ;
  		starting_line_per_granule:valid_min = -2147483648 ;
  		starting_line_per_granule:valid_max = 2147483647 ;
  		starting_line_per_granule:missing_value = -992, -993, -994, -995, -996, -997, -998, -999 ;
  		string starting_line_per_granule:long_name = "Index of the line that starts each granule" ;
  	double earthview_start_of_data(band, scans) ;
  		earthview_start_of_data:_FillValue = -999.8 ;
  		earthview_start_of_data:valid_min = 1.48323e+15 ;
  		earthview_start_of_data:valid_max = 2.27215e+15 ;
  		earthview_start_of_data:missing_value = -999.2, -999.3, -999.4, -999.5, -999.6, -999.7, -999.8, -999.9 ;
  		string earthview_start_of_data:coordinates = "band" ;
  		string earthview_start_of_data:units = "microseconds since 1958/01/01 00:00:00" ;
  		string earthview_start_of_data:long_name = "Time at scan start" ;
  		string earthview_start_of_data:source = "(APID805, APID809, APID807, APID808, APID810, APID812, APID816, APID815, APID814):TimeOfDayStartOfData" ;
  		string earthview_start_of_data:standard_name = "time" ;
  	double earthview_scan_terminus(band, scans) ;
  		earthview_scan_terminus:_FillValue = -999.8 ;
  		earthview_scan_terminus:valid_min = 1.48323e+15 ;
  		earthview_scan_terminus:valid_max = 2.27215e+15 ;
  		earthview_scan_terminus:missing_value = -999.2, -999.3, -999.4, -999.5, -999.6, -999.7, -999.8, -999.9 ;
  		string earthview_scan_terminus:coordinates = "band" ;
  		string earthview_scan_terminus:units = "microseconds since 1958/01/01 00:00:00" ;
  		string earthview_scan_terminus:long_name = "Time at scan terminus" ;
  		string earthview_scan_terminus:source = "(APID805, APID809, APID807, APID808, APID810, APID812, APID816, APID815, APID814):ScanTerminus" ;
  		string earthview_scan_terminus:standard_name = "time" ;
  	double calibview_start_of_data(calib_band, scans) ;
  		calibview_start_of_data:_FillValue = -999.8 ;
  		calibview_start_of_data:valid_min = 1.48323e+15 ;
  		calibview_start_of_data:valid_max = 2.27215e+15 ;
  		calibview_start_of_data:missing_value = -999.2, -999.3, -999.4, -999.5, -999.6, -999.7, -999.8, -999.9 ;
  		string calibview_start_of_data:coordinates = "calib_band" ;
  		string calibview_start_of_data:units = "microseconds since 1958/01/01 00:00:00" ;
  		string calibview_start_of_data:long_name = "Time at scan start" ;
  		string calibview_start_of_data:source = "APID825:TimeOfDayStartOfData (for each included band)" ;
  		string calibview_start_of_data:standard_name = "time" ;
  	double calibview_scan_terminus(calib_band, scans) ;
  		calibview_scan_terminus:_FillValue = -999.8 ;
  		calibview_scan_terminus:valid_min = 1.48323e+15 ;
  		calibview_scan_terminus:valid_max = 2.27215e+15 ;
  		calibview_scan_terminus:missing_value = -999.2, -999.3, -999.4, -999.5, -999.6, -999.7, -999.8, -999.9 ;
  		string calibview_scan_terminus:coordinates = "calib_band" ;
  		string calibview_scan_terminus:units = "microseconds since 1958/01/01 00:00:00" ;
  		string calibview_scan_terminus:long_name = "Time at scan terminus" ;
  		string calibview_scan_terminus:source = "APID825:ScanTerminus (for each included band)" ;
  		string calibview_scan_terminus:standard_name = "time" ;
  	uint earthview_band_control_word(band, scans) ;
  		earthview_band_control_word:_FillValue = 4294967294U ;
  		earthview_band_control_word:valid_min = 0U ;
  		earthview_band_control_word:valid_max = 4294967295U ;
  		earthview_band_control_word:missing_value = 4294967288U, 0U, 4294967289U, 0U, 4294967290U, 0U, 4294967291U, 0U ;
  		string earthview_band_control_word:coordinates = "band earthview_start_of_data" ;
  		string earthview_band_control_word:long_name = "Earth view Band Control Word" ;
  		string earthview_band_control_word:source = "(APID805, APID809, APID807, APID808, APID810, APID812, APID816, APID815, APID814):BandControlWord" ;
  	uint calibview_band_control_word(calib_band, scans) ;
  		calibview_band_control_word:_FillValue = 4294967294U ;
  		calibview_band_control_word:valid_min = 0U ;
  		calibview_band_control_word:valid_max = 4294967295U ;
  		calibview_band_control_word:missing_value = 4294967288U, 0U, 4294967289U, 0U, 4294967290U, 0U, 4294967291U, 0U ;
  		string calibview_band_control_word:coordinates = "calib_band calibview_start_of_data" ;
  		string calibview_band_control_word:long_name = "Calibration view Band Control Word" ;
  		string calibview_band_control_word:source = "APID825:BandControlWord (for each included band)" ;
  	ushort earthview(band, line, pixel) ;
  		earthview:_FillValue = 65534US ;
  		earthview:valid_min = 0US ;
  		earthview:valid_max = 4095US ;
  		earthview:missing_value = 65528US, 65529US, 65530US, 65531US, 65532US, 65533US, 65534US, 65535US ;
  		string earthview:coordinates = "band earthview_start_of_data" ;
  		string earthview:long_name = "Digital counts from the Earth view for Moderate single gain bands 6, 8-12, 14-16" ;
  		string earthview:source = "APID805, APID809, APID807, APID808, APID810, APID812, APID816, APID815, APID814" ;
  		earthview:chunk_size = 1, 3072, 3200 ;
  		earthview:chunk_compression_level = 2 ;
  	ushort calibview(calib_band, calib_source, line, cal_samples) ;
  		calibview:_FillValue = 65534US ;
  		calibview:valid_min = 0US ;
  		calibview:valid_max = 16383US ;
  		calibview:missing_value = 65528US, 65529US, 65530US, 65531US, 65532US, 65533US, 65534US, 65535US ;
  		string calibview:coordinates = "calib_band calib_source calibview_start_of_data" ;
  		string calibview:long_name = "Digital counts from the space view, black body, and solar diffuser for Moderate single gain bands 6, 8-12, 14-16" ;
  		string calibview:source = "APID825" ;
  		calibview:chunk_size = 1, 3, 3072, 48 ;
  		calibview:chunk_compression_level = 2 ;
  } // group Image_750m_SingleGain

group: Image_DayNight {
  dimensions:
  	line = UNLIMITED ; // (3072 currently)
  	pixel = 4064 ;
  	calib_source = 3 ;
  	cal_samples = 64 ;
  variables:
  	string calib_source(calib_source) ;
  		string calib_source:long_name = "calibration source identifier" ;
  	int lines_per_granule(granules) ;
  		lines_per_granule:_FillValue = -998 ;
  		lines_per_granule:valid_min = -2147483648 ;
  		lines_per_granule:valid_max = 2147483647 ;
  		lines_per_granule:missing_value = -992, -993, -994, -995, -996, -997, -998, -999 ;
  		string lines_per_granule:long_name = "Number of lines for each granule" ;
  	int starting_line_per_granule(granules) ;
  		starting_line_per_granule:_FillValue = -998 ;
  		starting_line_per_granule:valid_min = -2147483648 ;
  		starting_line_per_granule:valid_max = 2147483647 ;
  		starting_line_per_granule:missing_value = -992, -993, -994, -995, -996, -997, -998, -999 ;
  		string starting_line_per_granule:long_name = "Index of the line that starts each granule" ;
  	double earthview_start_of_data(scans) ;
  		earthview_start_of_data:_FillValue = -999.8 ;
  		earthview_start_of_data:valid_min = 1.48323e+15 ;
  		earthview_start_of_data:valid_max = 2.27215e+15 ;
  		earthview_start_of_data:missing_value = -999.2, -999.3, -999.4, -999.5, -999.6, -999.7, -999.8, -999.9 ;
  		string earthview_start_of_data:units = "microseconds since 1958/01/01 00:00:00" ;
  		string earthview_start_of_data:long_name = "Time at scan start" ;
  		string earthview_start_of_data:source = "APID821:TimeOfDayStartOfData" ;
  		string earthview_start_of_data:standard_name = "time" ;
  	double earthview_scan_terminus(scans) ;
  		earthview_scan_terminus:_FillValue = -999.8 ;
  		earthview_scan_terminus:valid_min = 1.48323e+15 ;
  		earthview_scan_terminus:valid_max = 2.27215e+15 ;
  		earthview_scan_terminus:missing_value = -999.2, -999.3, -999.4, -999.5, -999.6, -999.7, -999.8, -999.9 ;
  		string earthview_scan_terminus:units = "microseconds since 1958/01/01 00:00:00" ;
  		string earthview_scan_terminus:long_name = "Time at scan terminus" ;
  		string earthview_scan_terminus:source = "APID821:ScanTerminus" ;
  		string earthview_scan_terminus:standard_name = "time" ;
  	double calibview_start_of_data(scans) ;
  		calibview_start_of_data:_FillValue = -999.8 ;
  		calibview_start_of_data:valid_min = 1.48323e+15 ;
  		calibview_start_of_data:valid_max = 2.27215e+15 ;
  		calibview_start_of_data:missing_value = -999.2, -999.3, -999.4, -999.5, -999.6, -999.7, -999.8, -999.9 ;
  		string calibview_start_of_data:units = "microseconds since 1958/01/01 00:00:00" ;
  		string calibview_start_of_data:long_name = "Time at scan start" ;
  		string calibview_start_of_data:source = "APID825:TimeOfDayStartOfData (for Day/Night band)" ;
  		string calibview_start_of_data:standard_name = "time" ;
  	double calibview_scan_terminus(scans) ;
  		calibview_scan_terminus:_FillValue = -999.8 ;
  		calibview_scan_terminus:valid_min = 1.48323e+15 ;
  		calibview_scan_terminus:valid_max = 2.27215e+15 ;
  		calibview_scan_terminus:missing_value = -999.2, -999.3, -999.4, -999.5, -999.6, -999.7, -999.8, -999.9 ;
  		string calibview_scan_terminus:units = "microseconds since 1958/01/01 00:00:00" ;
  		string calibview_scan_terminus:long_name = "Time at scan terminus" ;
  		string calibview_scan_terminus:source = "APID825:ScanTerminus (for Day/Night band)" ;
  		string calibview_scan_terminus:standard_name = "time" ;
  	uint earthview_band_control_word(scans) ;
  		earthview_band_control_word:_FillValue = 4294967294U ;
  		earthview_band_control_word:valid_min = 0U ;
  		earthview_band_control_word:valid_max = 4294967295U ;
  		earthview_band_control_word:missing_value = 4294967288U, 0U, 4294967289U, 0U, 4294967290U, 0U, 4294967291U, 0U ;
  		string earthview_band_control_word:coordinates = "earthview_start_of_data" ;
  		string earthview_band_control_word:long_name = "Earth view Band Control Word" ;
  		string earthview_band_control_word:source = "APID821:BandControlWord" ;
  	uint calibview_band_control_word(scans) ;
  		calibview_band_control_word:_FillValue = 4294967294U ;
  		calibview_band_control_word:valid_min = 0U ;
  		calibview_band_control_word:valid_max = 4294967295U ;
  		calibview_band_control_word:missing_value = 4294967288U, 0U, 4294967289U, 0U, 4294967290U, 0U, 4294967291U, 0U ;
  		string calibview_band_control_word:coordinates = "calibview_start_of_data" ;
  		string calibview_band_control_word:long_name = "Calibration view Band Control Word" ;
  		string calibview_band_control_word:source = "APID825:BandControlWord (for Day/Night Band)" ;
  	ubyte calibview_dnb_agg_mode(scans) ;
  		calibview_dnb_agg_mode:_FillValue = 254UB ;
  		calibview_dnb_agg_mode:valid_min = 1UB ;
  		calibview_dnb_agg_mode:valid_max = 36UB ;
  		calibview_dnb_agg_mode:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string calibview_dnb_agg_mode:coordinates = "calibview_start_of_data" ;
  		string calibview_dnb_agg_mode:long_name = "Calibration Day/Night Band Aggregation Mode" ;
  		string calibview_dnb_agg_mode:source = "APID825:DNBAggMode" ;
  	ubyte calibview_active_samples(scans) ;
  		calibview_active_samples:_FillValue = 254UB ;
  		calibview_active_samples:valid_min = 0UB ;
  		calibview_active_samples:valid_max = 255UB ;
  		calibview_active_samples:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string calibview_active_samples:coordinates = "calibview_start_of_data" ;
  		string calibview_active_samples:long_name = "Active Day/Night Band calibration view samples per scan" ;
  	ushort earthview(line, pixel) ;
  		earthview:_FillValue = 65534US ;
  		earthview:valid_min = 0US ;
  		earthview:valid_max = 16383US ;
  		earthview:missing_value = 65528US, 65529US, 65530US, 65531US, 65532US, 65533US, 65534US, 65535US ;
  		string earthview:coordinates = "earthview_start_of_data" ;
  		string earthview:long_name = "Digital counts from the Earth view for Day/Night band" ;
  		string earthview:source = "APID821" ;
  		earthview:chunk_size = 3072, 4064 ;
  		earthview:chunk_compression_level = 2 ;
  	ubyte earthview_gain(line, pixel) ;
  		earthview_gain:_FillValue = 254UB ;
  		earthview_gain:valid_min = 0UB ;
  		earthview_gain:valid_max = 2UB ;
  		earthview_gain:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string earthview_gain:coordinates = "earthview_start_of_data" ;
  		string earthview_gain:long_name = "Gain state from the Earth view for Day/Night band" ;
  		string earthview_gain:source = "APID821" ;
  		earthview_gain:chunk_size = 3072, 4064 ;
  		earthview_gain:chunk_compression_level = 2 ;
  	ushort calibview(calib_source, line, cal_samples) ;
  		calibview:_FillValue = 65534US ;
  		calibview:valid_min = 0US ;
  		calibview:valid_max = 16383US ;
  		calibview:missing_value = 65528US, 65529US, 65530US, 65531US, 65532US, 65533US, 65534US, 65535US ;
  		string calibview:coordinates = "calib_source calibview_start_of_data" ;
  		string calibview:long_name = "Digital counts from the space view, black body, and solar diffuser for Day/Night band" ;
  		string calibview:source = "APID825" ;
  		calibview:chunk_size = 3, 3072, 64 ;
  		calibview:chunk_compression_level = 2 ;
  	ubyte calibview_gain(calib_source, line, cal_samples) ;
  		calibview_gain:_FillValue = 254UB ;
  		calibview_gain:valid_min = 0UB ;
  		calibview_gain:valid_max = 2UB ;
  		calibview_gain:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string calibview_gain:coordinates = "calib_source calibview_start_of_data" ;
  		string calibview_gain:long_name = "Gain state from the space view, black body, and solar diffuser for Day/Night band" ;
  		string calibview_gain:source = "APID825" ;
  		calibview_gain:chunk_size = 3, 3072, 64 ;
  		calibview_gain:chunk_compression_level = 2 ;
  } // group Image_DayNight

group: Quality_Measures {
  variables:
  	int scans_per_granule(granules) ;
  		scans_per_granule:_FillValue = -998 ;
  		scans_per_granule:valid_min = -2147483648 ;
  		scans_per_granule:valid_max = 2147483647 ;
  		scans_per_granule:missing_value = -992, -993, -994, -995, -996, -997, -998, -999 ;
  		string scans_per_granule:long_name = "Number of scans for each granule" ;
  	int starting_scan_per_granule(granules) ;
  		starting_scan_per_granule:_FillValue = -998 ;
  		starting_scan_per_granule:valid_min = -2147483648 ;
  		starting_scan_per_granule:valid_max = 2147483647 ;
  		starting_scan_per_granule:missing_value = -992, -993, -994, -995, -996, -997, -998, -999 ;
  		string starting_scan_per_granule:long_name = "Index of the scan that starts each granule" ;
  	int num_of_missing_packets(scans) ;
  		num_of_missing_packets:_FillValue = -998 ;
  		num_of_missing_packets:valid_min = 0 ;
  		num_of_missing_packets:valid_max = 2147483647 ;
  		num_of_missing_packets:missing_value = -992, -993, -994, -995, -996, -997, -998, -999 ;
  		string num_of_missing_packets:long_name = "Number of missing packets per scan" ;
  	int num_of_bad_checksums(scans) ;
  		num_of_bad_checksums:_FillValue = -998 ;
  		num_of_bad_checksums:valid_min = 0 ;
  		num_of_bad_checksums:valid_max = 2147483647 ;
  		num_of_bad_checksums:missing_value = -992, -993, -994, -995, -996, -997, -998, -999 ;
  		string num_of_bad_checksums:long_name = "Number of bad checksums per scan" ;
  	int num_of_discarded_packets(scans) ;
  		num_of_discarded_packets:_FillValue = -998 ;
  		num_of_discarded_packets:valid_min = 0 ;
  		num_of_discarded_packets:valid_max = 2147483647 ;
  		num_of_discarded_packets:missing_value = -992, -993, -994, -995, -996, -997, -998, -999 ;
  		string num_of_discarded_packets:long_name = "Number of discarded packets per scan" ;
  	uint rdr_scan_quality(scans) ;
  		rdr_scan_quality:_FillValue = 4294967294U ;
  		rdr_scan_quality:valid_min = 0U ;
  		rdr_scan_quality:valid_max = 4294967295U ;
  		rdr_scan_quality:missing_value = 4294967288U, 0U, 4294967289U, 0U, 4294967290U, 0U, 4294967291U, 0U ;
  		string rdr_scan_quality:long_name = "Quality flags for each scan" ;
  		rdr_scan_quality:flag_masks = 1, 2, 4, 8, 16, 32, 64 ;
  		string rdr_scan_quality:flag_meanings = "BadAggZone1 BadAggZone2 BadAggZone3 BadAggZone4 BadAggZone5 BadAggZone6 NoData" ;
  } // group Quality_Measures

group: Spacecraft_Diary {
  dimensions:
  	spacecraft_diary_granules = UNLIMITED ; // (18 currently)
  	bus_critical_sample = UNLIMITED ; // (360 currently)
  	adcs_hk_sample = UNLIMITED ; // (360 currently)
  	eph_att_sample = UNLIMITED ; // (360 currently)
  	ecf_axis = 3 ;
  	quaternion_element = 4 ;
  variables:
  	double bus_critical_packet_time(bus_critical_sample) ;
  		bus_critical_packet_time:_FillValue = -999.8 ;
  		bus_critical_packet_time:valid_min = 1.48323e+15 ;
  		bus_critical_packet_time:valid_max = 2.27215e+15 ;
  		bus_critical_packet_time:missing_value = -999.2, -999.3, -999.4, -999.5, -999.6, -999.7, -999.8, -999.9 ;
  		string bus_critical_packet_time:units = "microseconds since 1958/01/01 00:00:00" ;
  		string bus_critical_packet_time:long_name = "Bus Critical Telemetry packet time" ;
  		string bus_critical_packet_time:source = "APID0:TimeOfDayStartOfData" ;
  		string bus_critical_packet_time:standard_name = "time" ;
  	ubyte adcs_state(bus_critical_sample) ;
  		adcs_state:_FillValue = 254UB ;
  		adcs_state:valid_min = 0UB ;
  		adcs_state:valid_max = 4UB ;
  		adcs_state:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string adcs_state:coordinates = "bus_critical_packet_time" ;
  		string adcs_state:long_name = "Current ADCS State" ;
  		string adcs_state:source = "APID0:ADSTATE" ;
  		adcs_state:flag_values = 0b, 1b, 2b, 3b, 4b ;
  		string adcs_state:flag_meanings = "Wait/yel Detumble AcqSun Point DeltaV" ;
  	double adcs_hk_packet_time(adcs_hk_sample) ;
  		adcs_hk_packet_time:_FillValue = -999.8 ;
  		adcs_hk_packet_time:valid_min = 1.48323e+15 ;
  		adcs_hk_packet_time:valid_max = 2.27215e+15 ;
  		adcs_hk_packet_time:missing_value = -999.2, -999.3, -999.4, -999.5, -999.6, -999.7, -999.8, -999.9 ;
  		string adcs_hk_packet_time:units = "microseconds since 1958/01/01 00:00:00" ;
  		string adcs_hk_packet_time:long_name = "ADCS Housekeeping Telemetry packet time" ;
  		string adcs_hk_packet_time:source = "APID8:TimeOfDayStartOfData" ;
  		string adcs_hk_packet_time:standard_name = "time" ;
  	ubyte manuever_done(adcs_hk_sample) ;
  		manuever_done:_FillValue = 254UB ;
  		manuever_done:valid_min = 0UB ;
  		manuever_done:valid_max = 1UB ;
  		manuever_done:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
  		string manuever_done:coordinates = "adcs_hk_packet_time" ;
  		string manuever_done:long_name = "Maneuver Done state" ;
  		string manuever_done:source = "APID8:ADMANDONE" ;
  		manuever_done:flag_values = 0b, 1b ;
  		string manuever_done:flag_meanings = "Maneuver Done" ;
  	ushort fixed_frame_table_target_id(adcs_hk_sample) ;
  		fixed_frame_table_target_id:_FillValue = 65534US ;
  		fixed_frame_table_target_id:valid_min = 0US ;
  		fixed_frame_table_target_id:valid_max = 65535US ;
  		fixed_frame_table_target_id:missing_value = 65528US, 65529US, 65530US, 65531US, 65532US, 65533US, 65534US, 65535US ;
  		string fixed_frame_table_target_id:coordinates = "adcs_hk_packet_time" ;
  		string fixed_frame_table_target_id:long_name = "Fixed Frame Table Target ID" ;
  		string fixed_frame_table_target_id:source = "APID8:ADFFTID" ;
  	double ephemeris_valid_time(eph_att_sample) ;
  		ephemeris_valid_time:_FillValue = -999.8 ;
  		ephemeris_valid_time:valid_min = 1.48323e+15 ;
  		ephemeris_valid_time:valid_max = 2.27215e+15 ;
  		ephemeris_valid_time:missing_value = -999.2, -999.3, -999.4, -999.5, -999.6, -999.7, -999.8, -999.9 ;
  		string ephemeris_valid_time:units = "microseconds since 1958/01/01 00:00:00" ;
  		string ephemeris_valid_time:long_name = "ephemeris time" ;
  		string ephemeris_valid_time:source = "APID11:EphemerisValidTime" ;
  		string ephemeris_valid_time:standard_name = "time" ;
  	float ephemeris_position(eph_att_sample, ecf_axis) ;
  		ephemeris_position:_FillValue = -999.8f ;
  		ephemeris_position:valid_min = -7250000.f ;
  		ephemeris_position:valid_max = 7250000.f ;
  		ephemeris_position:missing_value = -999.2f, -999.3f, -999.4f, -999.5f, -999.6f, -999.7f, -999.8f, -999.9f ;
  		string ephemeris_position:coordinates = "ephemeris_valid_time" ;
  		string ephemeris_position:units = "meters" ;
  		string ephemeris_position:long_name = "Satellite position (ECEF)" ;
  		string ephemeris_position:source = "APID11:EphemerisPosition" ;
  	float ephemeris_velocity(eph_att_sample, ecf_axis) ;
  		ephemeris_velocity:_FillValue = -999.8f ;
  		ephemeris_velocity:valid_min = -7550.f ;
  		ephemeris_velocity:valid_max = 7550.f ;
  		ephemeris_velocity:missing_value = -999.2f, -999.3f, -999.4f, -999.5f, -999.6f, -999.7f, -999.8f, -999.9f ;
  		string ephemeris_velocity:coordinates = "ephemeris_valid_time" ;
  		string ephemeris_velocity:units = "m/s" ;
  		string ephemeris_velocity:long_name = "Satellite velocity (ECEF)" ;
  		string ephemeris_velocity:source = "APID11:EphemerisVelocity" ;
  	double attitude_valid_time(eph_att_sample) ;
  		attitude_valid_time:_FillValue = -999.8 ;
  		attitude_valid_time:valid_min = 1.48323e+15 ;
  		attitude_valid_time:valid_max = 2.27215e+15 ;
  		attitude_valid_time:missing_value = -999.2, -999.3, -999.4, -999.5, -999.6, -999.7, -999.8, -999.9 ;
  		string attitude_valid_time:units = "microseconds since 1958/01/01 00:00:00" ;
  		string attitude_valid_time:long_name = "attitude time" ;
  		string attitude_valid_time:source = "APID11:AttitudeValidTime" ;
  		string attitude_valid_time:standard_name = "time" ;
  	float control_frame_attitude_quaternion(eph_att_sample, quaternion_element) ;
  		control_frame_attitude_quaternion:_FillValue = -999.8f ;
  		control_frame_attitude_quaternion:valid_min = -1.f ;
  		control_frame_attitude_quaternion:valid_max = 1.f ;
  		control_frame_attitude_quaternion:missing_value = -999.2f, -999.3f, -999.4f, -999.5f, -999.6f, -999.7f, -999.8f, -999.9f ;
  		string control_frame_attitude_quaternion:coordinates = "attitude_valid_time" ;
  		string control_frame_attitude_quaternion:long_name = "Satellite orientation (ECI J2000.0)" ;
  		string control_frame_attitude_quaternion:source = "APID11:ControlFrameAttitudeQuaternions" ;

  // group attributes:
  		:Beginning_Orbit_Numbers = 23876U, 23876U, 23876U, 23876U, 23876U, 23876U, 23876U, 23876U, 23876U, 23876U, 23876U, 23876U, 23876U, 23876U, 23876U, 23876U, 23876U, 23876U ;
  		string :Input_RDR_Granule_IDs = "NPP001458688600", "NPP001458688800", "NPP001458689000", "NPP001458689200", "NPP001458689400", "NPP001458689600", "NPP001458689800", "NPP001458690000", "NPP001458690200", "NPP001458690400", "NPP001458690600", "NPP001458690800", "NPP001458691000", "NPP001458691200", "NPP001458691400", "NPP001458691600", "NPP001458691800", "NPP001458692000" ;
  		string :Input_RDR_Granule_Versions = "A1", "A1", "A1", "A1", "A1", "A1", "A1", "A1", "A1", "A1", "A1", "A1", "A1", "A1", "A1", "A1", "A1", "A1" ;
  		string :LEOA_Flags = "Off", "Off", "Off", "Off", "Off", "Off", "Off", "Off", "Off", "Off", "Off", "Off", "Off", "Off", "Off", "Off", "Off", "Off" ;
  		:Percent_Missing_Data = 4.7619f, 4.7619f, 4.7619f, 4.7619f, 4.7619f, 4.7619f, 4.7619f, 4.7619f, 4.7619f, 4.7619f, 4.7619f, 4.7619f, 4.7619f, 4.7619f, 4.7619f, 4.7619f, 4.7619f, 4.7619f ;

  group: ADCS_Housekeeping_Telemetry {
    dimensions:
    	packet_bytes = UNLIMITED ; // (355 currently)
    variables:
    	ubyte packets_per_granule(spacecraft_diary_granules) ;
    		packets_per_granule:_FillValue = 254UB ;
    		packets_per_granule:valid_min = 0UB ;
    		packets_per_granule:valid_max = 255UB ;
    		packets_per_granule:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
    		string packets_per_granule:long_name = "Number of ADCS Housekeeping Telemetry packets (APID 8) per Spacecraft Diary granule" ;
    		string packets_per_granule:source = "Spacecraft Diary RDR" ;
    	ushort starting_packet_per_granule(spacecraft_diary_granules) ;
    		starting_packet_per_granule:_FillValue = 65534US ;
    		starting_packet_per_granule:valid_min = 0US ;
    		starting_packet_per_granule:valid_max = 65535US ;
    		starting_packet_per_granule:missing_value = 65528US, 65529US, 65530US, 65531US, 65532US, 65533US, 65534US, 65535US ;
    		string starting_packet_per_granule:long_name = "Index of the first ADCS Housekeeping Telemetry packet for each Spacecraft Diary granule" ;
    	ushort packet_sequence_counter(adcs_hk_sample) ;
    		packet_sequence_counter:_FillValue = 65534US ;
    		packet_sequence_counter:valid_min = 0US ;
    		packet_sequence_counter:valid_max = 16383US ;
    		packet_sequence_counter:missing_value = 65528US, 65529US, 65530US, 65531US, 65532US, 65533US, 65534US, 65535US ;
    		string packet_sequence_counter:coordinates = "start_of_scan_time" ;
    		string packet_sequence_counter:long_name = "ADCS Housekeeping Telemetry Packet Sequence Count" ;
    		string packet_sequence_counter:source = "APID8:PacketSequenceCounter" ;
    	ubyte fill_percent(adcs_hk_sample) ;
    		fill_percent:_FillValue = 254UB ;
    		fill_percent:valid_min = 0UB ;
    		fill_percent:valid_max = 100UB ;
    		fill_percent:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
    		string fill_percent:coordinates = "packet_sequence_counter start_of_scan_time" ;
    		string fill_percent:units = "percent" ;
    		string fill_percent:long_name = "ADCS Housekeeping Telemetry fill percentage per packet" ;
    		string fill_percent:source = "Spacecraft Diary RDR" ;
    	ubyte packet(adcs_hk_sample, packet_bytes) ;
    		packet:_FillValue = 254UB ;
    		packet:valid_min = 0UB ;
    		packet:valid_max = 255UB ;
    		packet:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
    		string packet:coordinates = "packet_sequence_counter start_of_scan_time" ;
    		string packet:long_name = "ADCS Housekeeping Telemetry packet (APID 8)" ;
    		string packet:source = "APID8" ;
    } // group ADCS_Housekeeping_Telemetry

  group: Bus_Critical_Telemetry {
    dimensions:
    	packet_bytes = UNLIMITED ; // (207 currently)
    variables:
    	ubyte packets_per_granule(spacecraft_diary_granules) ;
    		packets_per_granule:_FillValue = 254UB ;
    		packets_per_granule:valid_min = 0UB ;
    		packets_per_granule:valid_max = 255UB ;
    		packets_per_granule:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
    		string packets_per_granule:long_name = "Number of Bus Critical Telemetry packets (APID 0) per Spacecraft Diary granule" ;
    		string packets_per_granule:source = "Spacecraft Diary RDR" ;
    	ushort starting_packet_per_granule(spacecraft_diary_granules) ;
    		starting_packet_per_granule:_FillValue = 65534US ;
    		starting_packet_per_granule:valid_min = 0US ;
    		starting_packet_per_granule:valid_max = 65535US ;
    		starting_packet_per_granule:missing_value = 65528US, 65529US, 65530US, 65531US, 65532US, 65533US, 65534US, 65535US ;
    		string starting_packet_per_granule:long_name = "Index of the first Bus Critical Telemetry packet for each Spacecraft Diary granule" ;
    	ushort packet_sequence_counter(bus_critical_sample) ;
    		packet_sequence_counter:_FillValue = 65534US ;
    		packet_sequence_counter:valid_min = 0US ;
    		packet_sequence_counter:valid_max = 16383US ;
    		packet_sequence_counter:missing_value = 65528US, 65529US, 65530US, 65531US, 65532US, 65533US, 65534US, 65535US ;
    		string packet_sequence_counter:coordinates = "packet_sequence_counter start_of_scan_time" ;
    		string packet_sequence_counter:long_name = "Bus Critical Telemetry Packet Sequence Count" ;
    		string packet_sequence_counter:source = "APID0:PacketSequenceCounter" ;
    	ubyte fill_percent(bus_critical_sample) ;
    		fill_percent:_FillValue = 254UB ;
    		fill_percent:valid_min = 0UB ;
    		fill_percent:valid_max = 100UB ;
    		fill_percent:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
    		string fill_percent:coordinates = "packet_sequence_counter start_of_scan_time" ;
    		string fill_percent:units = "percent" ;
    		string fill_percent:long_name = "Bus Critical Telemetry fill percentage per packet" ;
    		string fill_percent:source = "Spacecraft Diary RDR" ;
    	ubyte packet(bus_critical_sample, packet_bytes) ;
    		packet:_FillValue = 254UB ;
    		packet:valid_min = 0UB ;
    		packet:valid_max = 255UB ;
    		packet:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
    		string packet:coordinates = "packet_sequence_counter start_of_scan_time" ;
    		string packet:long_name = "Bus Critical Telemetry packet (APID 0)" ;
    		string packet:source = "APID0" ;
    } // group Bus_Critical_Telemetry

  group: Ephemeris_Attitude_Telemetry {
    dimensions:
    	packet_bytes = UNLIMITED ; // (71 currently)
    variables:
    	ubyte packets_per_granule(spacecraft_diary_granules) ;
    		packets_per_granule:_FillValue = 254UB ;
    		packets_per_granule:valid_min = 0UB ;
    		packets_per_granule:valid_max = 255UB ;
    		packets_per_granule:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
    		string packets_per_granule:long_name = "Number of Ephemeris/Attitude packets (APID 11) per Spacecraft Diary granule" ;
    		string packets_per_granule:source = "Spacecraft Diary RDR" ;
    	ushort starting_packet_per_granule(spacecraft_diary_granules) ;
    		starting_packet_per_granule:_FillValue = 65534US ;
    		starting_packet_per_granule:valid_min = 0US ;
    		starting_packet_per_granule:valid_max = 65535US ;
    		starting_packet_per_granule:missing_value = 65528US, 65529US, 65530US, 65531US, 65532US, 65533US, 65534US, 65535US ;
    		string starting_packet_per_granule:long_name = "Index of the first Ephemeris/Attitude packet for each Spacecraft Diary granule" ;
    	ushort packet_sequence_counter(eph_att_sample) ;
    		packet_sequence_counter:_FillValue = 65534US ;
    		packet_sequence_counter:valid_min = 0US ;
    		packet_sequence_counter:valid_max = 16383US ;
    		packet_sequence_counter:missing_value = 65528US, 65529US, 65530US, 65531US, 65532US, 65533US, 65534US, 65535US ;
    		string packet_sequence_counter:coordinates = "packet_sequence_counter start_of_scan_time" ;
    		string packet_sequence_counter:long_name = "Ephemeris/Attitude Packet Sequence Count" ;
    		string packet_sequence_counter:source = "APID11:PacketSequenceCounter" ;
    	ubyte fill_percent(eph_att_sample) ;
    		fill_percent:_FillValue = 254UB ;
    		fill_percent:valid_min = 0UB ;
    		fill_percent:valid_max = 100UB ;
    		fill_percent:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
    		string fill_percent:coordinates = "packet_sequence_counter start_of_scan_time" ;
    		string fill_percent:units = "percent" ;
    		string fill_percent:long_name = "Ephemeris/Attitude fill percentage per packet" ;
    		string fill_percent:source = "Spacecraft Diary RDR" ;
    	ubyte packet(eph_att_sample, packet_bytes) ;
    		packet:_FillValue = 254UB ;
    		packet:valid_min = 0UB ;
    		packet:valid_max = 255UB ;
    		packet:missing_value = 248UB, 249UB, 250UB, 251UB, 252UB, 253UB, 254UB, 255UB ;
    		string packet:coordinates = "packet_sequence_counter start_of_scan_time" ;
    		string packet:long_name = "Ephemeris/Attitude Telemetry packet (APID 11)" ;
    		string packet:source = "APID11" ;
    } // group Ephemeris_Attitude_Telemetry
  } // group Spacecraft_Diary
}
