netcdf S5P_TEST_L1B_RA_BD6_20140827T114200_20140827T115800_53811_01_000901_20141209T120000 {

		:time_coverage_end = "2014-08-27T11:51:47Z" ;
		:time_coverage_start = "2014-08-27T11:45:53Z" ;
		:time_reference = "2014-08-27T00:00:00Z" ;

group: BAND6_RADIANCE {

  group: STANDARD_MODE {
    dimensions:
    	time = 1 ;
    	scanline = 326 ; // flight direction
    	spectral_channel = 497 ; // spectral dimension
    	ground_pixel = 448 ; // scan direction (perpendicular to flight direction)
    	ncorner = 4 ;
    	nsettings = 5 ;
    	nbinningregions = 18 ;

    group: OBSERVATIONS {
      types:
        float(*) vlen_float ;
      variables:
      	int scanline(scanline) ;
      		scanline:comment = "This dimension variable defines the indices along track; index starts at 0" ;
      		scanline:long_name = "along track dimension index" ;
      		scanline:units = "1" ;
      	int delta_time(time, scanline) ;
      		delta_time:comment = "Time difference with time for each measurement" ;
      		delta_time:_FillValue = -2147483647 ;
      		delta_time:long_name = "offset from the reference start time of measurement" ;
      		delta_time:units = "milliseconds since 2014-08-27 00:00:00" ;
      	int spectral_channel(spectral_channel) ;
      		spectral_channel:comment = "This dimension variable defines the indices spectral dimension; index starts at 0" ;
      		spectral_channel:long_name = "wavelength dimension index" ;
      		spectral_channel:units = "1" ;
      	ushort detector_column_qualification(time, scanline, spectral_channel) ;
      		detector_column_qualification:comment = "Qualification flag indicating column indicating column type or state" ;
      		detector_column_qualification:units = "1" ;
      		detector_column_qualification:_FillValue = 65535US ;
      		detector_column_qualification:flag_values = 0US, 1US, 16US, 32US, 64US, 256US, 512US, 1024US, 2048US ;
      		detector_column_qualification:flag_masks = 0US, 1US, 16US, 98US, 98US, 3840US, 3840US, 3840US, 3840US ;
      		detector_column_qualification:flag_meanings = "no_qualification skipped uvn_odd uvn_prepost uvn_overscan swir_adc0 swir_adc1 swir_adc2 swir_adc3" ;
      		detector_column_qualification:long_name = "Detector column qualification flags" ;
      		detector_column_qualification:max_val = 65534US ;
      		detector_column_qualification:min_val = 0US ;
      	int ground_pixel(ground_pixel) ;
      		ground_pixel:comment = "This dimension variable defines the indices across track; index starts at 0" ;
      		ground_pixel:long_name = "across track dimension index" ;
      		ground_pixel:units = "1" ;
      	ushort detector_row_qualification(time, scanline, ground_pixel) ;
      		detector_row_qualification:comment = "Qualification flag indicating row type or state" ;
      		detector_row_qualification:_FillValue = 65535US ;
      		detector_row_qualification:flag_values = 0US, 1US, 2US, 4US, 8US, 16US, 256US, 4096US, 8192US ;
      		detector_row_qualification:flag_masks = 0US, 9US, 2US, 4US, 9US, 16US, 256US, 4096US, 8192US ;
      		detector_row_qualification:flag_meanings = "no_qualification uvn_ror uvn_dump uvn_covered uvn_overscan uvn_higain swir_reference gen_transistion gen_non_illuminated" ;
      		detector_row_qualification:long_name = "Detector row qualification flags" ;
      		detector_row_qualification:max_val = 65534US ;
      		detector_row_qualification:min_val = 0US ;
      		detector_row_qualification:units = "1" ;
      	ubyte ground_pixel_quality(time, scanline, ground_pixel) ;
      		ground_pixel_quality:comment = "Quality assessment information for each ground pixel" ;
      		ground_pixel_quality:coordinates = "longitude latitude" ;
      		ground_pixel_quality:max_val = 254UB ;
      		ground_pixel_quality:_FillValue = 255UB ;
      		ground_pixel_quality:flag_values = 0UB, 1UB, 2UB, 4UB, 8UB, 16UB, 128UB ;
      		ground_pixel_quality:flag_masks = 0UB, 1UB, 2UB, 4UB, 8UB, 16UB, 128UB ;
      		ground_pixel_quality:flag_meanings = "no_error solar_eclipse sun_glint_possible descending night geo_boundary_crossing geolocation_error" ;
      		ground_pixel_quality:long_name = "ground pixel quality flag" ;
      		ground_pixel_quality:min_val = 0UB ;
      		ground_pixel_quality:units = "1" ;
      	ushort measurement_quality(time, scanline) ;
      		measurement_quality:flag_masks = 0US, 1US, 2US, 16US, 32US, 128US, 256US, 4096US ;
      		measurement_quality:flag_meanings = "no_error proc_skipped no_residual saa spacecraft_manoeuvre sub_grp irr_out_of_range sub_group" ;
      		measurement_quality:long_name = "measurement quality flag" ;
      		measurement_quality:max_val = 65534US ;
      		measurement_quality:min_val = 0US ;
      		measurement_quality:units = "1" ;
      		measurement_quality:comment = "Overall quality information for a measurement" ;
      		measurement_quality:coordinates = "longitude latitude" ;
      		measurement_quality:_FillValue = 65535US ;
      		measurement_quality:flag_values = 0US, 1US, 2US, 16US, 32US, 128US, 256US, 4096US ;
      	ubyte quality_level(time, scanline, ground_pixel, spectral_channel) ;
      		quality_level:comment = "Overall quality assessment information for each (spectral) pixel" ;
      		quality_level:coordinates = "longitude latitude" ;
      		quality_level:_FillValue = 255UB ;
      		quality_level:long_name = "qualiy level of spectral channel" ;
      		quality_level:max_val = 100UB ;
      		quality_level:min_val = 0UB ;
      		quality_level:units = "1" ;
      	float radiance(time, scanline, ground_pixel, spectral_channel) ;
      		radiance:ancilary_vars = "radiance_noise radiance_error quality_level spectral_channel_quality ground_pixel_quality" ;
      		radiance:coordinates = "longitude latitude" ;
      		radiance:comment = "Measured spectral radiance for each spectral pixel" ;
      		radiance:_FillValue = 9.96921e+36f ;
      		radiance:long_name = "spectral photon radiance" ;
      		radiance:units = "mol.m-2.nm-1.sr-1.s-1" ;
      	byte radiance_error(time, scanline, ground_pixel, spectral_channel) ;
      		radiance_error:comment = "The radiance_error is a measure for the one standard deviation error of the bias of the radiance measurement; it is expressed in decibel (dB), i.e. 10 times the base-10 logarithmic value of the ratio between the radiance and the estimation error." ;
      		radiance_error:coordinates = "longitude latitude" ;
      		radiance_error:_FillValue = -127b ;
      		radiance_error:long_name = "spectral photon radiance error, one standard deviation" ;
      		radiance_error:units = "1" ;
      	byte radiance_noise(time, scanline, ground_pixel, spectral_channel) ;
      		radiance_noise:coordinates = "longitude latitude" ;
      		radiance_noise:comment = "The radiance_noise is a measure for the one standard deviation random error of the radiance measurement; it is expressed in decibel (dB), i.e. 10 times the base-10 logarithmic value of the ratio between the radiance and the random error." ;
      		radiance_noise:_FillValue = -127b ;
      		radiance_noise:long_name = "spectral photon radiance noise, one standard deviation" ;
      		radiance_noise:units = "1" ;
      	vlen_float small_pixel_radiance(time, scanline, ground_pixel) ;
      		small_pixel_radiance:long_name = "small pixel photon radiance" ;
      		small_pixel_radiance:units = "mol.m-2.nm-1.sr-1.s-1" ;
      		small_pixel_radiance:comment = "Measured spectral radiance for the spectral channel dedicated for the small pixel measurements" ;
      		small_pixel_radiance:coordinates = "longitude latitude" ;
      	ubyte spectral_channel_quality(time, scanline, ground_pixel, spectral_channel) ;
      		spectral_channel_quality:comment = "Quality assessment information for each (spectral) pixel" ;
      		spectral_channel_quality:units = "1" ;
      		spectral_channel_quality:coordinates = "longitude latitude" ;
      		spectral_channel_quality:_FillValue = 255UB ;
      		spectral_channel_quality:flag_values = 0UB, 1UB, 2UB, 8UB, 16UB, 32UB, 64UB, 128UB ;
      		spectral_channel_quality:flag_masks = 0UB, 1UB, 2UB, 8UB, 16UB, 32UB, 64UB, 128UB ;
      		spectral_channel_quality:flag_meanings = "no_error missing bad_pixel processing_error saturated transient rts underflow" ;
      		spectral_channel_quality:long_name = "spectral channel quality flag" ;
      		spectral_channel_quality:max_val = 254UB ;
      		spectral_channel_quality:min_val = 0UB ;
      	int time(time) ;
      		time:comment = "Reference time of the measurements. The reference time is set to yyyy-mm-ddT00:00:00 UTC, where yyyy-mm-dd is the day on which the measurements of a particular data granule start." ;
      		time:long_name = "reference start time of measurement" ;
      		time:standard_name = "time" ;
      		time:units = "seconds since 2010-01-01 00:00:00" ;
      } // group OBSERVATIONS

    group: GEODATA {
      variables:
      	float earth_sun_distance(time) ;
      		earth_sun_distance:comment = "1 ua equals 149,597,870,700 meters" ;
      		earth_sun_distance:_FillValue = 9.96921e+36f ;
      		earth_sun_distance:units = "ua" ;
      		earth_sun_distance:long_name = "distance between the earth and the sun" ;
      		earth_sun_distance:max_val = 1.02f ;
      		earth_sun_distance:min_val = 0.98f ;
      	float latitude_bounds(time, scanline, ground_pixel, ncorner) ;
      		latitude_bounds:comment = "The four latitude boundaries of each ground pixel." ;
      		latitude_bounds:_FillValue = 9.96921e+36f ;
      		latitude_bounds:units = "degrees north" ;
      	float latitude(time, scanline, ground_pixel) ;
      		latitude:comment = "Latitude of the center of each ground pixel on the WGS84  reference ellipsoid" ;
      		latitude:_FillValue = 9.96921e+36f ;
      		latitude:long_name = "pixel center latitude" ;
      		latitude:max_val = 90.f ;
      		latitude:min_val = -90.f ;
      		latitude:standard_name = "latitude" ;
      		latitude:bounds = "latitude_bounds" ;
      		latitude:units = "degrees north" ;
      	float longitude_bounds(time, scanline, ground_pixel, ncorner) ;
      		longitude_bounds:comment = "The four longitude boundaries of each ground pixel." ;
      		longitude_bounds:_FillValue = 9.96921e+36f ;
      		longitude_bounds:units = "degrees east" ;
      	float longitude(time, scanline, ground_pixel) ;
      		longitude:comment = "Longitude of the center of each ground pixel on the WGS84 reference ellipsoid" ;
      		longitude:_FillValue = 9.96921e+36f ;
      		longitude:long_name = "pixel center longitude" ;
      		longitude:bounds = "longitude_bounds" ;
      		longitude:max_val = 180.f ;
      		longitude:min_val = -180.f ;
      		longitude:standard_name = "longitude" ;
      		longitude:units = "degrees east" ;
      	float satellite_altitude(time, scanline) ;
      		satellite_altitude:comment = "The altitude of the spacecraft relative to the WGS84 reference ellipsoid" ;
      		satellite_altitude:_FillValue = 9.96921e+36f ;
      		satellite_altitude:long_name = "satellite altitude" ;
      		satellite_altitude:max_val = 900000.f ;
      		satellite_altitude:min_val = 700000.f ;
      		satellite_altitude:units = "m" ;
      	float satellite_latitude(time, scanline) ;
      		satellite_latitude:comment = "Latitude of the spacecraft sub-satellite point on the WGS84 reference ellipsoid" ;
      		satellite_latitude:_FillValue = 9.96921e+36f ;
      		satellite_latitude:long_name = "sub-satellite latitude" ;
      		satellite_latitude:max_val = 90.f ;
      		satellite_latitude:min_val = -90.f ;
      		satellite_latitude:units = "degrees north" ;
      	float satellite_longitude(time, scanline) ;
      		satellite_longitude:comment = "Longitude of the spacecraft sub-satellite point on the WGS84 reference ellipsoid" ;
      		satellite_longitude:_FillValue = 9.96921e+36f ;
      		satellite_longitude:max_val = 180.f ;
      		satellite_longitude:min_val = -180.f ;
      		satellite_longitude:units = "degrees east" ;
      	float satellite_orbit_phase(time, scanline) ;
      		satellite_orbit_phase:comment = "Relative offset (0.0 ... 1.0) of the measurement in the orbit" ;
      		satellite_orbit_phase:_FillValue = 9.96921e+36f ;
      		satellite_orbit_phase:long_name = "fractional satellite orbit phase" ;
      		satellite_orbit_phase:max_val = 1.02f ;
      		satellite_orbit_phase:min_val = -0.02f ;
      		satellite_orbit_phase:units = "1" ;
      	float solar_azimuth_angle(time, scanline, ground_pixel) ;
      		solar_azimuth_angle:units = "degree" ;
      		solar_azimuth_angle:comment = "Solar azimuth angle at the ground pixel location on the reference ellipsoid. Angle is measured clockwise from the North (East = 90, South = 180, West = 270)" ;
      		solar_azimuth_angle:coordinates = "longitude latitude" ;
      		solar_azimuth_angle:_FillValue = 9.96921e+36f ;
      		solar_azimuth_angle:long_name = "solar azimuth angle" ;
      		solar_azimuth_angle:max_val = 360.f ;
      		solar_azimuth_angle:min_val = 0.f ;
      		solar_azimuth_angle:standard_name = "solar_azimuth_angle" ;
      	float solar_zenith_angle(time, scanline, ground_pixel) ;
      		solar_zenith_angle:comment = "Solar zenith angle at the ground pixel location on the reference ellipsoid. Angle is measured away from the vertical. ESA definition of day side: SZA less the 92 degrees" ;
      		solar_zenith_angle:coordinates = "longitude latitude" ;
      		solar_zenith_angle:_FillValue = 9.96921e+36f ;
      		solar_zenith_angle:long_name = "solar zenith angle" ;
      		solar_zenith_angle:max_val = 180.f ;
      		solar_zenith_angle:min_val = 0.f ;
      		solar_zenith_angle:standard_name = "solar_zenith_angle" ;
      		solar_zenith_angle:units = "degree" ;
      	float viewing_azimuth_angle(time, scanline, ground_pixel) ;
      		viewing_azimuth_angle:comment = "Azimuth angle of the satellite at the ground pixel location on the reference ellipsoid. Angle is measured clockwise from the North (East = 90, South = 180, West = 270)" ;
      		viewing_azimuth_angle:coordinates = "longitude latitude" ;
      		viewing_azimuth_angle:_FillValue = 9.96921e+36f ;
      		viewing_azimuth_angle:units = "degree" ;
      		viewing_azimuth_angle:long_name = "viewing azimuth angle" ;
      		viewing_azimuth_angle:max_val = 360.f ;
      		viewing_azimuth_angle:min_val = 0.f ;
      		viewing_azimuth_angle:standard_name = "platform_azimuth_angle" ;
      	float viewing_zenith_angle(time, scanline, ground_pixel) ;
      		viewing_zenith_angle:comment = "Zenith angle of the satellite at the ground pixel location on the reference ellipsoid. Angle is measured away from the vertical." ;
      		viewing_zenith_angle:coordinates = "longitude latitude" ;
      		viewing_zenith_angle:_FillValue = 9.96921e+36f ;
      		viewing_zenith_angle:long_name = "viewing zenith angle" ;
      		viewing_zenith_angle:max_val = 180.f ;
      		viewing_zenith_angle:min_val = 0.f ;
      		viewing_zenith_angle:standard_name = "platform_zenith_angle" ;
      		viewing_zenith_angle:units = "degree" ;
      } // group GEODATA

    } // group STANDARD_MODE
  } // group BAND6_RADIANCE
}
