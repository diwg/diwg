// Contributed by Jessica Hausman <Jessica.K.Hausman AT jpl DOT nasa DOT gov>

netcdf Q2015005015300 {

// global attributes:
		:Product\ Name = "Q2015005015300.L1A_SCI" ;
		:Title = "Aquarius Level 1A Data" ;
		:Data\ Center = "NASA/GSFC Aquarius Data Processing Center" ;
		:Mission = "SAC-D Aquarius" ;
		:Mission\ Characteristics = "Nominal orbit: inclination=98.0 (Sun-synchronous); node=6PM (ascending); eccentricity=<0.002; altitude=657 km; ground speed=6.825 km/sec" ;
		:Sensor = "Aquarius" ;
		:Data\ Type = "SCI" ;
		:Software\ ID = "1.05" ;
		:Processing\ Time = "2015006124942000" ;
		:Input\ Files = "Q20150105_095106_T20150105_000500_20150105_020259.AQ_L1A,Q20150105_095106_T20150105_014301_20150105_034058.AQ_L1A,Q20150105_095106_T20150105_032100_20150105_051859.AQ_L1A,Q20150105_043731_T20150105_000500_20150105_020259.AQ_L1A,Q20150105_043731_T20150105_014301_20150105_034058.AQ_L1A,Q20150105_043731_T20150105_032100_20150105_043731.AQ_L1A" ;
		:Processing\ Control = "l1amerge_aquarius l1amerge.inputs /data7/sdpsoper/vdc/vpu6/workbuf" ;
		:Number\ of\ Beams = 3 ;
		:Radiometer\ Polarizations = 4 ;
		:Radiometer\ Subcycles = 12 ;
		:Radiometer\ Signals\ per\ Subcycle = 5 ;
		:Radiometer\ Long\ Accumulations = 8 ;
		:Scatterometer\ Polarizations = 6 ;
		:Scatterometer\ Subcycles = 8 ;
		:Start\ Time = "2015005014301309" ;
		:Start\ Year = 2015 ;
		:Start\ Day = 5 ;
		:Start\ Millisec = 6181309 ;
		:End\ Year = 2015 ;
		:End\ Day = 5 ;
		:End\ Millisec = 13258911 ;
		:Orbit\ Start\ Time = "2015005015300000" ;
		:Orbit\ Stop\ Time = "2015005033100000" ;
		:Number\ of\ Orbit\ Vectors = 120 ;
		:Number\ of\ Attitude\ Samples = 887 ;
		:Number\ of\ Blocks = 4916 ;
		:Number\ of\ RAD\ Frames = 1229 ;
		:Number\ of\ ATC\ Frames = 1229 ;
		:End\ Time = "2015005034058911" ;
		:Product\ Center\ Time = "2015005024200110" ;
		:Node\ Crossing\ Time = "2015005021730000" ;
		:Orbit\ Number = 19195 ;
		:Cycle\ Number = 176 ;
		:Pass\ Number = 61 ;
		:Orbit\ Node\ Longitude = -123.1856f ;
		:Radiometer\ LUTs\ Block\ Count = 4916, 0, 0, 0, 0, 0, 0, 0 ;
		:Percent\ Non-default\ Radiometer\ LUTs = 0.f ;
		:Missing\ Blocks = 0 ;

group: Block\ Attributes {
  dimensions:
  	phony_dim_0 = 5200 ;
  variables:
  	int atc_frmnum(phony_dim_0) ;
  		atc_frmnum:long_name = "ATC Frame Number" ;
  		atc_frmnum:valid_min = 0 ;
  		atc_frmnum:valid_max = 0 ;
  	ubyte atc_subframe(phony_dim_0) ;
  		atc_subframe:long_name = "ATC Sub-Frame Number" ;
  		atc_subframe:valid_min = 0UB ;
  		atc_subframe:valid_max = 0UB ;
  	double blk_sec(phony_dim_0) ;
  		blk_sec:long_name = "Block time, seconds of day" ;
  		blk_sec:valid_min = 0. ;
  		blk_sec:valid_max = 0. ;
  		blk_sec:units = "seconds" ;
  	int rad_frmnum(phony_dim_0) ;
  		rad_frmnum:long_name = "Radiometer Frame Number" ;
  		rad_frmnum:valid_min = 0 ;
  		rad_frmnum:valid_max = 0 ;
  	ubyte rad_subframe(phony_dim_0) ;
  		rad_subframe:long_name = "Radiometer Sub-Frame Number" ;
  		rad_subframe:valid_max = 0UB ;
  		rad_subframe:valid_min = 0UB ;
  } // group Block\ Attributes

group: Converted\ Telemetry {
  dimensions:
  	phony_dim_1 = 5200 ;
  	phony_dim_2 = 5 ;
  	phony_dim_3 = 1300 ;
  	phony_dim_4 = 17 ;
  	phony_dim_5 = 4 ;
  	phony_dim_6 = 7 ;
  	phony_dim_7 = 12 ;
  	phony_dim_8 = 13 ;
  	phony_dim_9 = 38 ;
  	phony_dim_10 = 14 ;
  	phony_dim_11 = 8 ;
  	phony_dim_12 = 21 ;
  	phony_dim_13 = 23 ;
  	phony_dim_14 = 30 ;
  variables:
  	float apdu_analog_tlm(phony_dim_1, phony_dim_2) ;
  		apdu_analog_tlm:long_name = "Aquarius Power Distribution Unit analog telemetry" ;
  		apdu_analog_tlm:valid_min = 0.f ;
  		apdu_analog_tlm:valid_max = 0.f ;
  	float atc_omt1_analog_tlm(phony_dim_3, phony_dim_4) ;
  		atc_omt1_analog_tlm:long_name = "ATC OMT1 analog telemetry" ;
  		atc_omt1_analog_tlm:valid_min = 0.f ;
  		atc_omt1_analog_tlm:valid_max = 0.f ;
  	ubyte atc_omt1_discrete_tlm(phony_dim_3, phony_dim_4) ;
  		atc_omt1_discrete_tlm:long_name = "ATC OMT1 discrete telemetry" ;
  		atc_omt1_discrete_tlm:valid_min = 0UB ;
  		atc_omt1_discrete_tlm:valid_max = 0UB ;
  	float atc_omt2_analog_tlm(phony_dim_3, phony_dim_4) ;
  		atc_omt2_analog_tlm:long_name = "ATC OMT2 analog telemetry" ;
  		atc_omt2_analog_tlm:valid_min = 0.f ;
  		atc_omt2_analog_tlm:valid_max = 0.f ;
  	ubyte atc_omt2_discrete_tlm(phony_dim_3, phony_dim_4) ;
  		atc_omt2_discrete_tlm:long_name = "ATC OMT2 discrete telemetry" ;
  		atc_omt2_discrete_tlm:valid_min = 0UB ;
  		atc_omt2_discrete_tlm:valid_max = 0UB ;
  	float atc_omt3_analog_tlm(phony_dim_3, phony_dim_4) ;
  		atc_omt3_analog_tlm:long_name = "ATC OMT3 analog telemetry" ;
  		atc_omt3_analog_tlm:valid_min = 0.f ;
  		atc_omt3_analog_tlm:valid_max = 0.f ;
  	ubyte atc_omt3_discrete_tlm(phony_dim_3, phony_dim_4) ;
  		atc_omt3_discrete_tlm:long_name = "ATC OMT3 discrete telemetry" ;
  		atc_omt3_discrete_tlm:valid_min = 0UB ;
  		atc_omt3_discrete_tlm:valid_max = 0UB ;
  	float atc_rbe_analog_tlm(phony_dim_3, phony_dim_4) ;
  		atc_rbe_analog_tlm:long_name = "ATC RBE analog telemetry" ;
  		atc_rbe_analog_tlm:valid_min = 0.f ;
  		atc_rbe_analog_tlm:valid_max = 0.f ;
  	ubyte atc_rbe_discrete_tlm(phony_dim_3, phony_dim_4) ;
  		atc_rbe_discrete_tlm:long_name = "ATC RBE discrete telemetry" ;
  		atc_rbe_discrete_tlm:valid_min = 0UB ;
  		atc_rbe_discrete_tlm:valid_max = 0UB ;
  	float deploy_analog_tlm(phony_dim_1, phony_dim_5) ;
  		deploy_analog_tlm:long_name = "Antenna deployment analog telemetry" ;
  		deploy_analog_tlm:valid_min = 0.f ;
  		deploy_analog_tlm:valid_max = 0.f ;
  	int deploy_discrete_tlm(phony_dim_1, phony_dim_6) ;
  		deploy_discrete_tlm:long_name = "Antenna deployment discrete telemetry" ;
  		deploy_discrete_tlm:valid_min = 0 ;
  		deploy_discrete_tlm:valid_max = 0 ;
  	float dpu_analog_tlm(phony_dim_3, phony_dim_7) ;
  		dpu_analog_tlm:long_name = "DPU analog telemetry" ;
  		dpu_analog_tlm:valid_min = 0.f ;
  		dpu_analog_tlm:valid_max = 0.f ;
  	ubyte dpu_status_tlm(phony_dim_3, phony_dim_5, phony_dim_8) ;
  		dpu_status_tlm:long_name = "DPU discrete telemetry" ;
  		dpu_status_tlm:valid_min = 0UB ;
  		dpu_status_tlm:valid_max = 0UB ;
  	float ext_temp_analog_tlm(phony_dim_1, phony_dim_9) ;
  		ext_temp_analog_tlm:long_name = "External Temperature Sensor analog telemetry" ;
  		ext_temp_analog_tlm:valid_min = 0.f ;
  		ext_temp_analog_tlm:valid_max = 0.f ;
  	float icds_analog_tlm(phony_dim_1, phony_dim_10) ;
  		icds_analog_tlm:long_name = "ICDS analog telemetry" ;
  		icds_analog_tlm:valid_max = 0.f ;
  		icds_analog_tlm:valid_min = 0.f ;
  	int icds_discrete_tlm(phony_dim_1, phony_dim_11) ;
  		icds_discrete_tlm:long_name = "ICDS discrete telemetry" ;
  		icds_discrete_tlm:valid_min = 0 ;
  		icds_discrete_tlm:valid_max = 0 ;
  	ushort radiom_nrt_tlm(phony_dim_3, phony_dim_5, phony_dim_4) ;
  		radiom_nrt_tlm:long_name = "Radiometer discrete non-real-time telemetry" ;
  		radiom_nrt_tlm:valid_min = 0US ;
  		radiom_nrt_tlm:valid_max = 0US ;
  	float rbe1_analog_tlm(phony_dim_3, phony_dim_12) ;
  		rbe1_analog_tlm:long_name = "RBE1 analog telemetry" ;
  		rbe1_analog_tlm:valid_min = 0.f ;
  		rbe1_analog_tlm:valid_max = 0.f ;
  	float rbe2_analog_tlm(phony_dim_3, phony_dim_12) ;
  		rbe2_analog_tlm:long_name = "RBE2 analog telemetry" ;
  		rbe2_analog_tlm:valid_min = 0.f ;
  		rbe2_analog_tlm:valid_max = 0.f ;
  	float rbe3_analog_tlm(phony_dim_3, phony_dim_12) ;
  		rbe3_analog_tlm:long_name = "RBE3 analog telemetry" ;
  		rbe3_analog_tlm:valid_max = 0.f ;
  		rbe3_analog_tlm:valid_min = 0.f ;
  	float rfe1_analog_tlm(phony_dim_3, phony_dim_13) ;
  		rfe1_analog_tlm:long_name = "RFE1 analog telemetry" ;
  		rfe1_analog_tlm:valid_max = 0.f ;
  		rfe1_analog_tlm:valid_min = 0.f ;
  	float rfe2_analog_tlm(phony_dim_3, phony_dim_13) ;
  		rfe2_analog_tlm:long_name = "RFE2 analog telemetry" ;
  		rfe2_analog_tlm:valid_min = 0.f ;
  		rfe2_analog_tlm:valid_max = 0.f ;
  	float rfe3_analog_tlm(phony_dim_3, phony_dim_13) ;
  		rfe3_analog_tlm:long_name = "RFE3 analog telemetry" ;
  		rfe3_analog_tlm:valid_min = 0.f ;
  		rfe3_analog_tlm:valid_max = 0.f ;
  	float scatter_analog_tlm(phony_dim_1, phony_dim_14) ;
  		scatter_analog_tlm:long_name = "Scatterometer analog telemetry" ;
  		scatter_analog_tlm:valid_min = 0.f ;
  		scatter_analog_tlm:valid_max = 0.f ;
  	ubyte scatter_discrete_tlm(phony_dim_1, phony_dim_11) ;
  		scatter_discrete_tlm:long_name = "Scatterometer discrete telemetry" ;
  		scatter_discrete_tlm:valid_max = 0UB ;
  		scatter_discrete_tlm:valid_min = 0UB ;
  } // group Converted\ Telemetry

group: Navigation {
  dimensions:
  	phony_dim_15 = 937 ;
  	phony_dim_16 = 3 ;
  	phony_dim_17 = 125 ;
  	phony_dim_18 = 4 ;
  variables:
  	double att_ang(phony_dim_15, phony_dim_16) ;
  		att_ang:long_name = "Spacecraft roll, pitch, yaw" ;
  		att_ang:valid_min = -180. ;
  		att_ang:valid_max = 180. ;
  		att_ang:units = "degrees" ;
  	int att_flags(phony_dim_15) ;
  		att_flags:long_name = "Attitude flags" ;
  		att_flags:valid_min = 0 ;
  		att_flags:valid_max = 0 ;
  	double att_time(phony_dim_15) ;
  		att_time:long_name = "Time tag of attitude data" ;
  		att_time:valid_min = 0. ;
  		att_time:valid_max = 0. ;
  		att_time:units = "seconds" ;
  	double orb_pos(phony_dim_17, phony_dim_16) ;
  		orb_pos:long_name = "Orbital position vector" ;
  		orb_pos:valid_min = -7100000. ;
  		orb_pos:valid_max = 7100000. ;
  		orb_pos:units = "meters" ;
  	double orb_time(phony_dim_17) ;
  		orb_time:long_name = "Time tag of orbit vectors" ;
  		orb_time:valid_min = 0. ;
  		orb_time:valid_max = 0. ;
  		orb_time:units = "seconds" ;
  	double orb_vel(phony_dim_17, phony_dim_16) ;
  		orb_vel:long_name = "Orbital velocity vector" ;
  		orb_vel:valid_min = -7600. ;
  		orb_vel:valid_max = 7600. ;
  		orb_vel:units = "meters per second" ;
  	double quaternion(phony_dim_15, phony_dim_18) ;
  		quaternion:long_name = "ECI-to-spacecraft quaternion" ;
  		quaternion:valid_max = 1. ;
  		quaternion:valid_min = -1. ;
  } // group Navigation

group: Raw\ Aquarius\ Data {
  dimensions:
  	phony_dim_19 = 5200 ;
  	phony_dim_20 = 5 ;
  	phony_dim_21 = 36 ;
  	phony_dim_22 = 12 ;
  	phony_dim_23 = 24 ;
  	phony_dim_24 = 35 ;
  	phony_dim_25 = 1300 ;
  	phony_dim_26 = 4 ;
  	phony_dim_27 = 3 ;
  	phony_dim_28 = 8 ;
  	phony_dim_29 = 10 ;
  	phony_dim_30 = 50 ;
  	phony_dim_31 = 2 ;
  	phony_dim_32 = 6 ;
  	phony_dim_33 = 37 ;
  	phony_dim_34 = 70 ;
  variables:
  	ubyte apdu_tlm(phony_dim_19, phony_dim_20) ;
  		apdu_tlm:long_name = "Aquarius Power Distribution Unit telemetry" ;
  		apdu_tlm:valid_min = 0UB ;
  		apdu_tlm:valid_max = 0UB ;
  	ubyte atc_tlm(phony_dim_19, phony_dim_21) ;
  		atc_tlm:long_name = "Active Thermal Control Unit telemetry" ;
  		atc_tlm:valid_min = 0UB ;
  		atc_tlm:valid_max = 0UB ;
  	ushort checksum(phony_dim_19) ;
  		checksum:long_name = "Checksum" ;
  		checksum:valid_min = 0US ;
  		checksum:valid_max = 0US ;
  	ubyte deploy_tlm(phony_dim_19, phony_dim_20) ;
  		deploy_tlm:long_name = "Antenna deployment telemetry" ;
  		deploy_tlm:valid_min = 0UB ;
  		deploy_tlm:valid_max = 0UB ;
  	int gps_time_tag(phony_dim_19) ;
  		gps_time_tag:long_name = "Block GPS time tag" ;
  		gps_time_tag:valid_min = 0 ;
  		gps_time_tag:valid_max = 0 ;
  		gps_time_tag:units = "seconds" ;
  	ubyte icds_status(phony_dim_19, phony_dim_22) ;
  		icds_status:long_name = "ICDS processing status" ;
  		icds_status:valid_min = 0UB ;
  		icds_status:valid_max = 0UB ;
  	ubyte icds_tlm(phony_dim_19, phony_dim_23) ;
  		icds_tlm:long_name = "ICDS engineering telemetry" ;
  		icds_tlm:valid_min = 0UB ;
  		icds_tlm:valid_max = 0UB ;
  	ubyte pad(phony_dim_19, phony_dim_24) ;
  		pad:long_name = "Pad" ;
  		pad:valid_min = 0UB ;
  		pad:valid_max = 0UB ;
  	ushort radiom_cnd(phony_dim_25, phony_dim_26, phony_dim_22, phony_dim_27, phony_dim_26) ;
  		radiom_cnd:long_name = "Radiometer CND Looks" ;
  		radiom_cnd:valid_min = 0US ;
  		radiom_cnd:valid_max = 0US ;
  	ushort radiom_header(phony_dim_25, phony_dim_26) ;
  		radiom_header:long_name = "Radiometer block header" ;
  		radiom_header:valid_min = 0US ;
  		radiom_header:valid_max = 0US ;
  	ushort radiom_lavg(phony_dim_25, phony_dim_26, phony_dim_28, phony_dim_27, phony_dim_26) ;
  		radiom_lavg:long_name = "Radiometer Long Accumulations" ;
  		radiom_lavg:valid_min = 0US ;
  		radiom_lavg:valid_max = 0US ;
  	ubyte radiom_nrt_tlm(phony_dim_25, phony_dim_26, phony_dim_29) ;
  		radiom_nrt_tlm:long_name = "Radiometer non-real-time telemetry" ;
  		radiom_nrt_tlm:valid_min = 0UB ;
  		radiom_nrt_tlm:valid_max = 0UB ;
  	ubyte radiom_rt_tlm(phony_dim_25, phony_dim_26, phony_dim_30) ;
  		radiom_rt_tlm:long_name = "Radiometer real-time telemetry" ;
  		radiom_rt_tlm:valid_min = 0UB ;
  		radiom_rt_tlm:valid_max = 0UB ;
  	ushort radiom_signals(phony_dim_25, phony_dim_26, phony_dim_22, phony_dim_20, phony_dim_27, phony_dim_26) ;
  		radiom_signals:long_name = "Radiometer Antenna Looks" ;
  		radiom_signals:valid_min = 0US ;
  		radiom_signals:valid_max = 0US ;
  	ushort scatter_dc(phony_dim_19, phony_dim_31) ;
  		scatter_dc:long_name = "Scatterometer DC data" ;
  		scatter_dc:valid_min = 0US ;
  		scatter_dc:valid_max = 0US ;
  	ubyte scatter_headers(phony_dim_19, phony_dim_28) ;
  		scatter_headers:long_name = "Scatterometer subcycle headers" ;
  		scatter_headers:valid_min = 0UB ;
  		scatter_headers:valid_max = 0UB ;
  	ushort scatter_loop(phony_dim_19, phony_dim_27, phony_dim_32) ;
  		scatter_loop:long_name = "Scatterometer Loopback Measurements" ;
  		scatter_loop:valid_min = 0US ;
  		scatter_loop:valid_max = 0US ;
  	ushort scatter_pwr(phony_dim_19, phony_dim_28, phony_dim_27, phony_dim_32) ;
  		scatter_pwr:long_name = "Scatterometer Power" ;
  		scatter_pwr:valid_min = 0US ;
  		scatter_pwr:valid_max = 0US ;
  	ubyte scatter_rfi(phony_dim_19, phony_dim_26) ;
  		scatter_rfi:long_name = "Scatterometer RFI flags for H-pol" ;
  		scatter_rfi:valid_min = 0UB ;
  		scatter_rfi:valid_max = 0UB ;
  	ubyte scatter_tlm(phony_dim_19, phony_dim_33) ;
  		scatter_tlm:long_name = "Scatterometer telemetry" ;
  		scatter_tlm:valid_min = 0UB ;
  		scatter_tlm:valid_max = 0UB ;
  	int start_synch(phony_dim_19) ;
  		start_synch:long_name = "Start-synch word" ;
  		start_synch:valid_min = 0 ;
  		start_synch:valid_max = 0 ;
  		start_synch:units = "dummy" ;
  	ubyte temp_tlm(phony_dim_19, phony_dim_34) ;
  		temp_tlm:long_name = "External Temperature Sensors telemetry" ;
  		temp_tlm:valid_min = 0UB ;
  		temp_tlm:valid_max = 0UB ;
  	int time_tag_offset(phony_dim_19) ;
  		time_tag_offset:long_name = "Block time offset from GPS" ;
  		time_tag_offset:valid_min = 0 ;
  		time_tag_offset:valid_max = 0 ;
  		time_tag_offset:units = "62.5 nanosec units" ;
  } // group Raw\ Aquarius\ Data

group: SAC-D\ Telemetry {
  dimensions:
  	phony_dim_35 = 1040 ;
  	phony_dim_36 = 4000 ;
  variables:
  	ubyte sacd_hkt(phony_dim_35, phony_dim_36) ;
  		sacd_hkt:long_name = "SAC-D raw housekeeping telemetry blocks" ;
  		sacd_hkt:valid_min = 0UB ;
  		sacd_hkt:valid_max = 0UB ;
  } // group SAC-D\ Telemetry
}
