// Contributed by Jessica Hausman <Jessica.K.Hausman AT jpl DOT nasa DOT gov>

netcdf JA1_GPN_2PeP073_013_20031230_143922_20031230_153534 {
dimensions:
	time = 3124 ;
	meas_ind = 20 ;
variables:
	double time(time) ;
		time:long_name = "time (sec. since 2000-01-01)" ;
		time:standard_name = "time" ;
		time:calendar = "gregorian" ;
		time:tai_utc_difference = 32. ;
		time:leap_second = "0000-00-00 00:00:00" ;
		time:units = "seconds since 2000-01-01 00:00:00.0" ;
		time:comment = "[tai_utc_difference] is the difference between TAI - UTC (i.e., leap seconds) for the first measurement of the data set. [leap_second] is the UTC time at which a leap second occurs in the data set, if any. After this UTC time, the [tai_utc_difference] is increased by 1 second. time variable is corrected from datation bias. See Jason-1 User handbook." ;
	byte meas_ind(meas_ind) ;
		meas_ind:long_name = "elementary measurement index" ;
		meas_ind:units = "count" ;
		meas_ind:comment = "Set to be compliant with the CF-1.1 convention" ;
	double time_20hz(time, meas_ind) ;
		time_20hz:_FillValue = 1.84467440737096e+19 ;
		time_20hz:long_name = "time 20 Hz (sec. since 2000-01-01)" ;
		time_20hz:standard_name = "time" ;
		time_20hz:calendar = "gregorian" ;
		time_20hz:tai_utc_difference = 32. ;
		time_20hz:leap_second = "0000-00-00 00:00:00" ;
		time_20hz:units = "seconds since 2000-01-01 00:00:00.0" ;
		time_20hz:comment = "[tai_utc_difference] is the difference between TAI - UTC (i.e., leap seconds) for the first measurement of the data set. [leap_second] is the UTC time at which a leap second occurs in the data set, if any. After this UTC time, the [tai_utc_difference] is increased by 1 second. time_20hz variable is corrected from datation bias. See Jason-1 User handbook." ;
	int lat(time) ;
		lat:long_name = "latitude" ;
		lat:standard_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:quality_flag = "orb_state_flag_rest" ;
		lat:scale_factor = 1.e-06 ;
		lat:comment = "Positive latitude is North latitude, negative latitude is South latitude. See Jason-1 User Handbook." ;
	int lon(time) ;
		lon:long_name = "longitude" ;
		lon:standard_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:quality_flag = "orb_state_flag_rest" ;
		lon:scale_factor = 1.e-06 ;
		lon:comment = "East longitude relative to Greenwich meridian. See Jason-1 User Handbook." ;
	int lon_20hz(time, meas_ind) ;
		lon_20hz:_FillValue = 2147483647 ;
		lon_20hz:long_name = "20 Hz longitude" ;
		lon_20hz:standard_name = "longitude" ;
		lon_20hz:units = "degrees_east" ;
		lon_20hz:scale_factor = 1.e-06 ;
		lon_20hz:comment = "East longitude relative to Greenwich meridian. See Jason-1 User Handbook" ;
	int lat_20hz(time, meas_ind) ;
		lat_20hz:_FillValue = 2147483647 ;
		lat_20hz:long_name = "20 Hz latitude" ;
		lat_20hz:standard_name = "latitude" ;
		lat_20hz:units = "degrees_north" ;
		lat_20hz:scale_factor = 1.e-06 ;
		lat_20hz:comment = "Positive latitude is North latitude, negative latitude is South latitude. See Jason-1 User Handbook" ;
	byte surface_type(time) ;
		surface_type:_FillValue = 127b ;
		surface_type:long_name = "surface type" ;
		surface_type:flag_values = 0b, 1b, 2b, 3b ;
		surface_type:flag_meanings = "ocean lake_enclosed_sea ice land" ;
		surface_type:coordinates = "lon lat" ;
		surface_type:comment = "Computed using a DTM2000 file: 0 = open oceans or semi-enclosed seas; 1 = enclosed seas or lakes; 2 = continental ice; 3 = land. See Jason-1 User Handbook" ;
	byte surface_type_globcover(time) ;
		surface_type_globcover:_FillValue = 127b ;
		surface_type_globcover:long_name = "surface type globcover" ;
		surface_type_globcover:flag_values = "0b, 1b, 2b, 3b, 4b, 5b, 6b" ;
		surface_type_globcover:flag_meanings = "open_ocean land continental_water aquatic_vegetation continental_ice_snow floating_ice salted_basin" ;
		surface_type_globcover:coordinates = "lon lat" ;
		surface_type_globcover:comment = "Computed from a mask built with MODIS and GlobCover data, 0 = Open ocean; 1 = Land; 2 = Continental waters; 3 = Aquatic vegetation; 4 = Continental ice and snow; 5 = Floating ice; 6 = Salted basin. See Jason-1 User Handbook" ;
	byte alt_echo_type(time) ;
		alt_echo_type:_FillValue = 127b ;
		alt_echo_type:long_name = "altimeter echo type" ;
		alt_echo_type:flag_values = 0b, 1b ;
		alt_echo_type:flag_meanings = "ocean_like non_ocean_like" ;
		alt_echo_type:coordinates = "lon lat" ;
		alt_echo_type:comment = "The altimeter echo type is determined by testing the rms of the high rate range measurements against a threshold as well as the number of valid high rate range measurements against a minimum value" ;
	byte rad_surf_type(time) ;
		rad_surf_type:_FillValue = 127b ;
		rad_surf_type:long_name = "radiometer surface type" ;
		rad_surf_type:flag_values = 0b, 1b, 2b ;
		rad_surf_type:flag_meanings = "open_ocean near_coast land" ;
		rad_surf_type:coordinates = "lon lat" ;
		rad_surf_type:comment = " The radiometer surface type flag is applicable to the radiometer wet troposphere path delays provided by rad_wet_tropo_corr. A value of 0 indicates that open ocean processing is used to compute the path delay, 1 indicates coastal processing is used, and 2 indicates the path delay is invalid due to land" ;
	int rad_distance_to_land(time) ;
		rad_distance_to_land:_FillValue = 2147483647 ;
		rad_distance_to_land:long_name = "radiometer radial distance to land" ;
		rad_distance_to_land:units = "m" ;
		rad_distance_to_land:coordinates = "lon lat" ;
		rad_distance_to_land:comment = "Shortest distance between nadir sub-satellite point and land" ;
	byte qual_alt_1hz_range_ku(time) ;
		qual_alt_1hz_range_ku:_FillValue = 127b ;
		qual_alt_1hz_range_ku:long_name = "quality flag for 1 Hz altimeter data: Ku band range" ;
		qual_alt_1hz_range_ku:flag_values = 0b, 1b ;
		qual_alt_1hz_range_ku:flag_meanings = "good bad" ;
		qual_alt_1hz_range_ku:coordinates = "lon lat" ;
	byte qual_alt_1hz_range_c(time) ;
		qual_alt_1hz_range_c:_FillValue = 127b ;
		qual_alt_1hz_range_c:long_name = "quality flag for 1 Hz altimeter data: C band range" ;
		qual_alt_1hz_range_c:flag_values = 0b, 1b ;
		qual_alt_1hz_range_c:flag_meanings = "good bad" ;
		qual_alt_1hz_range_c:coordinates = "lon lat" ;
	byte qual_alt_1hz_swh_ku(time) ;
		qual_alt_1hz_swh_ku:_FillValue = 127b ;
		qual_alt_1hz_swh_ku:long_name = "quality flag for 1 Hz altimeter data: Ku band SWH" ;
		qual_alt_1hz_swh_ku:flag_values = 0b, 1b ;
		qual_alt_1hz_swh_ku:flag_meanings = "good bad" ;
		qual_alt_1hz_swh_ku:coordinates = "lon lat" ;
	byte qual_alt_1hz_swh_c(time) ;
		qual_alt_1hz_swh_c:_FillValue = 127b ;
		qual_alt_1hz_swh_c:long_name = "quality flag for 1 Hz altimeter data: C band SWH" ;
		qual_alt_1hz_swh_c:flag_values = 0b, 1b ;
		qual_alt_1hz_swh_c:flag_meanings = "good bad" ;
		qual_alt_1hz_swh_c:coordinates = "lon lat" ;
	byte qual_alt_1hz_sig0_ku(time) ;
		qual_alt_1hz_sig0_ku:_FillValue = 127b ;
		qual_alt_1hz_sig0_ku:long_name = "quality flag for 1 Hz altimeter data: Ku band backscatter coefficient" ;
		qual_alt_1hz_sig0_ku:flag_values = 0b, 1b ;
		qual_alt_1hz_sig0_ku:flag_meanings = "good bad" ;
		qual_alt_1hz_sig0_ku:coordinates = "lon lat" ;
	byte qual_alt_1hz_sig0_c(time) ;
		qual_alt_1hz_sig0_c:_FillValue = 127b ;
		qual_alt_1hz_sig0_c:long_name = "quality flag for 1 Hz altimeter data: C band backscatter coefficient" ;
		qual_alt_1hz_sig0_c:flag_values = 0b, 1b ;
		qual_alt_1hz_sig0_c:flag_meanings = "good bad" ;
		qual_alt_1hz_sig0_c:coordinates = "lon lat" ;
	byte qual_alt_1hz_off_nadir_angle_wf_ku(time) ;
		qual_alt_1hz_off_nadir_angle_wf_ku:_FillValue = 127b ;
		qual_alt_1hz_off_nadir_angle_wf_ku:long_name = "quality flag for 1 Hz altimeter data: off nadir angle from Ku band" ;
		qual_alt_1hz_off_nadir_angle_wf_ku:flag_values = 0b, 1b ;
		qual_alt_1hz_off_nadir_angle_wf_ku:flag_meanings = "good bad" ;
		qual_alt_1hz_off_nadir_angle_wf_ku:coordinates = "lon lat" ;
	byte qual_inst_corr_1hz_range_ku(time) ;
		qual_inst_corr_1hz_range_ku:_FillValue = 127b ;
		qual_inst_corr_1hz_range_ku:long_name = "quality flag for 1 Hz instrumental correction: Ku band range" ;
		qual_inst_corr_1hz_range_ku:flag_values = 0b, 1b ;
		qual_inst_corr_1hz_range_ku:flag_meanings = "good bad" ;
		qual_inst_corr_1hz_range_ku:coordinates = "lon lat" ;
	byte qual_inst_corr_1hz_range_c(time) ;
		qual_inst_corr_1hz_range_c:_FillValue = 127b ;
		qual_inst_corr_1hz_range_c:long_name = "quality flag for 1 Hz instrumental correction: C band range" ;
		qual_inst_corr_1hz_range_c:flag_values = 0b, 1b ;
		qual_inst_corr_1hz_range_c:flag_meanings = "good bad" ;
		qual_inst_corr_1hz_range_c:coordinates = "lon lat" ;
	byte qual_inst_corr_1hz_swh_ku(time) ;
		qual_inst_corr_1hz_swh_ku:_FillValue = 127b ;
		qual_inst_corr_1hz_swh_ku:long_name = "quality flag for 1 Hz instrumental correction: Ku band SWH" ;
		qual_inst_corr_1hz_swh_ku:flag_values = 0b, 1b ;
		qual_inst_corr_1hz_swh_ku:flag_meanings = "good bad" ;
		qual_inst_corr_1hz_swh_ku:coordinates = "lon lat" ;
	byte qual_inst_corr_1hz_swh_c(time) ;
		qual_inst_corr_1hz_swh_c:_FillValue = 127b ;
		qual_inst_corr_1hz_swh_c:long_name = "quality flag for 1 Hz instrumental correction: C band SWH" ;
		qual_inst_corr_1hz_swh_c:flag_values = 0b, 1b ;
		qual_inst_corr_1hz_swh_c:flag_meanings = "good bad" ;
		qual_inst_corr_1hz_swh_c:coordinates = "lon lat" ;
	byte qual_inst_corr_1hz_sig0_ku(time) ;
		qual_inst_corr_1hz_sig0_ku:_FillValue = 127b ;
		qual_inst_corr_1hz_sig0_ku:long_name = "quality flag for 1 Hz instrumental correction: Ku band backscatter coefficient" ;
		qual_inst_corr_1hz_sig0_ku:flag_values = 0b, 1b ;
		qual_inst_corr_1hz_sig0_ku:flag_meanings = "good bad" ;
		qual_inst_corr_1hz_sig0_ku:coordinates = "lon lat" ;
	byte qual_inst_corr_1hz_sig0_c(time) ;
		qual_inst_corr_1hz_sig0_c:_FillValue = 127b ;
		qual_inst_corr_1hz_sig0_c:long_name = "quality flag for 1 Hz instrumental correction: C band backscatter coefficient" ;
		qual_inst_corr_1hz_sig0_c:flag_values = 0b, 1b ;
		qual_inst_corr_1hz_sig0_c:flag_meanings = "good bad" ;
		qual_inst_corr_1hz_sig0_c:coordinates = "lon lat" ;
	byte qual_rad_1hz_tb187(time) ;
		qual_rad_1hz_tb187:_FillValue = 127b ;
		qual_rad_1hz_tb187:long_name = "quality flag for 1 Hz radiometer data: 18.7 GHz brightness temperature" ;
		qual_rad_1hz_tb187:flag_values = 0b, 1b ;
		qual_rad_1hz_tb187:flag_meanings = "good bad" ;
		qual_rad_1hz_tb187:coordinates = "lon lat" ;
	byte qual_rad_1hz_tb238(time) ;
		qual_rad_1hz_tb238:_FillValue = 127b ;
		qual_rad_1hz_tb238:long_name = "quality flag for 1 Hz radiometer data: 23.8 GHz brightness temperature" ;
		qual_rad_1hz_tb238:flag_values = 0b, 1b ;
		qual_rad_1hz_tb238:flag_meanings = "good bad" ;
		qual_rad_1hz_tb238:coordinates = "lon lat" ;
	byte qual_rad_1hz_tb340(time) ;
		qual_rad_1hz_tb340:_FillValue = 127b ;
		qual_rad_1hz_tb340:long_name = "quality flag for 1 Hz radiometer data: 34.0 GHz brightness temperature" ;
		qual_rad_1hz_tb340:flag_values = 0b, 1b ;
		qual_rad_1hz_tb340:flag_meanings = "good bad" ;
		qual_rad_1hz_tb340:coordinates = "lon lat" ;
	byte rad_averaging_flag(time) ;
		rad_averaging_flag:_FillValue = 127b ;
		rad_averaging_flag:long_name = "radiometer along-track averaging flag" ;
		rad_averaging_flag:flag_values = 0b, 1b ;
		rad_averaging_flag:flag_meanings = "good bad" ;
		rad_averaging_flag:coordinates = "lon lat" ;
	short rad_land_frac_187(time) ;
		rad_land_frac_187:_FillValue = 32767s ;
		rad_land_frac_187:long_name = "radiometer 18.7 GHz antenna gain weighted land fraction in main beam" ;
		rad_land_frac_187:units = "%" ;
		rad_land_frac_187:scale_factor = 0.01 ;
		rad_land_frac_187:coordinates = "lon lat" ;
	short rad_land_frac_238(time) ;
		rad_land_frac_238:_FillValue = 32767s ;
		rad_land_frac_238:long_name = "radiometer 23.8 GHz antenna gain weighted land fraction in main beam" ;
		rad_land_frac_238:units = "%" ;
		rad_land_frac_238:scale_factor = 0.01 ;
		rad_land_frac_238:coordinates = "lon lat" ;
	short rad_land_frac_340(time) ;
		rad_land_frac_340:_FillValue = 32767s ;
		rad_land_frac_340:long_name = "radiometer 34.0 GHz antenna gain weighted land fraction in main beam" ;
		rad_land_frac_340:units = "%" ;
		rad_land_frac_340:scale_factor = 0.01 ;
		rad_land_frac_340:coordinates = "lon lat" ;
	byte alt_state_flag_oper(time) ;
		alt_state_flag_oper:_FillValue = 127b ;
		alt_state_flag_oper:long_name = "altimeter state flag: altimeter operating" ;
		alt_state_flag_oper:flag_values = 0b, 1b ;
		alt_state_flag_oper:flag_meanings = "SideA SideB" ;
		alt_state_flag_oper:coordinates = "lon lat" ;
		alt_state_flag_oper:comment = "Side A = nominal; Side B = redondancy" ;
	byte alt_state_flag_c_band(time) ;
		alt_state_flag_c_band:_FillValue = 127b ;
		alt_state_flag_c_band:long_name = "altimeter state flag: C bandwidth used" ;
		alt_state_flag_c_band:flag_values = 0b, 1b ;
		alt_state_flag_c_band:flag_meanings = "320MHz 100MHz" ;
		alt_state_flag_c_band:coordinates = "lon lat" ;
	byte alt_state_flag_band_seq(time) ;
		alt_state_flag_band_seq:_FillValue = 127b ;
		alt_state_flag_band_seq:long_name = "altimeter state flag: Ku/C band sequencing" ;
		alt_state_flag_band_seq:flag_values = 0b, 1b ;
		alt_state_flag_band_seq:flag_meanings = "3Ku_1C_3Ku 2Ku_1C_2Ku" ;
		alt_state_flag_band_seq:coordinates = "lon lat" ;
	byte alt_state_flag_ku_band_status(time) ;
		alt_state_flag_ku_band_status:_FillValue = 127b ;
		alt_state_flag_ku_band_status:long_name = "altimeter state flag: Ku band status" ;
		alt_state_flag_ku_band_status:flag_values = 0b, 1b ;
		alt_state_flag_ku_band_status:flag_meanings = "On Off" ;
		alt_state_flag_ku_band_status:coordinates = "lon lat" ;
	byte alt_state_flag_c_band_status(time) ;
		alt_state_flag_c_band_status:_FillValue = 127b ;
		alt_state_flag_c_band_status:long_name = "altimeter state flag: C band status" ;
		alt_state_flag_c_band_status:flag_values = 0b, 1b ;
		alt_state_flag_c_band_status:flag_meanings = "On Off" ;
		alt_state_flag_c_band_status:coordinates = "lon lat" ;
	byte rad_state_flag_oper(time) ;
		rad_state_flag_oper:_FillValue = 127b ;
		rad_state_flag_oper:long_name = "radiometer state flag: radiometer operating" ;
		rad_state_flag_oper:flag_values = 0b, 1b ;
		rad_state_flag_oper:flag_meanings = "Side A Side B" ;
		rad_state_flag_oper:coordinates = "lon lat" ;
		rad_state_flag_oper:comment = "Side A  nominal; Side B  redundancy" ;
	byte orb_state_flag_rest(time) ;
		orb_state_flag_rest:_FillValue = 127b ;
		orb_state_flag_rest:long_name = "orbit state flag: restituted orbit" ;
		orb_state_flag_rest:flag_values = 0b, 1b, 2b, 3b, 4b, 5b, 6b, 7b, 8b, 9b ;
		orb_state_flag_rest:flag_meanings = "op_maneuver op_adjusted op_extrapolated pre_adjusted pre_maneuver pre_interpolated_gap pre_extrapolated_L1 pre_extrapolated_L1S2 pre_extrapolated_S2 DIODE" ;
		orb_state_flag_rest:coordinates = "lon lat" ;
		orb_state_flag_rest:comment = "0 characterizes a mission operations orbit that is computed during a maneuver period, 1 stands for an adjusted mission operations orbit, 2 stands for an extrapolated mission operations orbit, 3 stands for an adjusted (preliminary/precise) orbit, 4 indicates that the (preliminary/precise) orbit is estimated during a maneuver period, 5 indicates that the (preliminary/precise) orbit is interpolated over a tracking data gap, 6 means that the (preliminary/precise) orbit is extrapolated for a duration less than 1 day, 7 means that the (preliminary/precise) orbit is extrapolated for a duration that ranges from 1 day to 2 days, 8 means that the (preliminary/precise) orbit is extrapolated for a duration larger than 2 days, or that the orbit is extrapolated just after a maneuver, 9 stands for the DORIS DIODE navigator orbit. The nominal value is 3" ;
	byte rain_flag(time) ;
		rain_flag:_FillValue = 127b ;
		rain_flag:long_name = "rain flag" ;
		rain_flag:flag_values = 0b, 1b ;
		rain_flag:flag_meanings = "no_rain rain" ;
		rain_flag:coordinates = "lon lat" ;
		rain_flag:comment = "See Jason-1 User Handbook" ;
	byte rad_rain_flag(time) ;
		rad_rain_flag:_FillValue = 127b ;
		rad_rain_flag:long_name = "radiometer rain flag" ;
		rad_rain_flag:flag_values = 0b, 1b ;
		rad_rain_flag:flag_meanings = "no_rain rain" ;
		rad_rain_flag:coordinates = "lon lat" ;
		rad_rain_flag:comment = "See Jason-1 User Handbook. The radiometer rain flag indicates where the radiometer wet troposphere path delay (rad_wet_tropo_corr) is invalid due to rain contamination" ;
	byte ice_flag(time) ;
		ice_flag:_FillValue = 127b ;
		ice_flag:long_name = "ice flag" ;
		ice_flag:flag_values = 0b, 1b ;
		ice_flag:flag_meanings = "no_ice ice" ;
		ice_flag:coordinates = "lon lat" ;
		ice_flag:comment = "See Jason-1 User Handbook" ;
	byte rad_sea_ice_flag(time) ;
		rad_sea_ice_flag:_FillValue = 127b ;
		rad_sea_ice_flag:long_name = "radiometer sea-ice flag" ;
		rad_sea_ice_flag:flag_values = 0b, 1b ;
		rad_sea_ice_flag:flag_meanings = "no_sea_ice, sea_ice" ;
		rad_sea_ice_flag:coordinates = "lon lat" ;
		rad_sea_ice_flag:comment = "See Jason-1 User Handbook. The radiometer sea ice flag indicates where the radiometer wet troposphere path delay (rad_wet_tropo_corr) is invalid due to sea ice contamination" ;
	byte interp_flag_tb(time) ;
		interp_flag_tb:_FillValue = 127b ;
		interp_flag_tb:long_name = "radiometer brightness temperatures interpolation flag" ;
		interp_flag_tb:flag_values = 0b, 1b, 2b, 3b ;
		interp_flag_tb:flag_meanings = "good interpolation_with_gap extrapolation fail" ;
		interp_flag_tb:coordinates = "lon lat" ;
		interp_flag_tb:comment = "Possible values are: 0  interpolation without gap between JMR data, 1 interpolation with gap between JMR data, 2  extrapolation of JMR data, 3  failure of extrapolation and interpolation" ;
	byte interp_flag_ocean_tide_sol1(time) ;
		interp_flag_ocean_tide_sol1:_FillValue = 127b ;
		interp_flag_ocean_tide_sol1:long_name = "ocean tide solution 1 interpolation flag" ;
		interp_flag_ocean_tide_sol1:flag_values = "0b, 1b" ;
		interp_flag_ocean_tide_sol1:flag_meanings = "good bad" ;
		interp_flag_ocean_tide_sol1:coordinates = "lon lat" ;
		interp_flag_ocean_tide_sol1:comment = "0 = valid interpolation; 1 = failure of interpolation i.e. ocean_tide_sol1 set to default value" ;
	byte interp_flag_ocean_tide_sol2(time) ;
		interp_flag_ocean_tide_sol2:_FillValue = 127b ;
		interp_flag_ocean_tide_sol2:long_name = "ocean tide solution 2 interpolation flag" ;
		interp_flag_ocean_tide_sol2:flag_values = "0b, 1b" ;
		interp_flag_ocean_tide_sol2:flag_meanings = "good bad" ;
		interp_flag_ocean_tide_sol2:coordinates = "lon lat" ;
		interp_flag_ocean_tide_sol2:comment = "0 = valid interpolation; 1 = failure of interpolation i.e. ocean_tide_sol2 set to default value" ;
	int alt(time) ;
		alt:_FillValue = 2147483647 ;
		alt:long_name = "1 Hz altitude of satellite" ;
		alt:standard_name = "height_above_reference_ellipsoid" ;
		alt:units = "m" ;
		alt:quality_flag = "orb_state_flag_rest" ;
		alt:add_offset = 1300000. ;
		alt:scale_factor = 0.0001 ;
		alt:coordinates = "lon lat" ;
		alt:comment = "Altitude of satellite above the reference ellipsoid." ;
	int alt_20hz(time, meas_ind) ;
		alt_20hz:_FillValue = 2147483647 ;
		alt_20hz:long_name = "20 Hz altitude of satellite" ;
		alt_20hz:standard_name = "height_above_reference_ellipsoid" ;
		alt_20hz:units = "m" ;
		alt_20hz:add_offset = 1300000. ;
		alt_20hz:scale_factor = 0.0001 ;
		alt_20hz:coordinates = "lon_20hz lat_20hz" ;
		alt_20hz:comment = "Altitude of satellite above reference ellipsoid" ;
	short orb_alt_rate(time) ;
		orb_alt_rate:_FillValue = 32767s ;
		orb_alt_rate:long_name = "1 Hz orbital altitude rate" ;
		orb_alt_rate:units = "m/s" ;
		orb_alt_rate:scale_factor = 0.01 ;
		orb_alt_rate:coordinates = "lon lat" ;
		orb_alt_rate:comment = "The reference surface for the orbital altitude rate is the combined mean_sea_surface/geoid surface. It is used to compute the Doppler correction on the altimeter range (doppler_corr_ku, doppler_corr_c)" ;
	int range_ku(time) ;
		range_ku:_FillValue = 2147483647 ;
		range_ku:long_name = "1 Hz Ku band corrected altimeter range" ;
		range_ku:standard_name = "altimeter_range" ;
		range_ku:units = "m" ;
		range_ku:quality_flag = "qual_alt_1hz_range_ku" ;
		range_ku:add_offset = 1300000. ;
		range_ku:scale_factor = 0.0001 ;
		range_ku:coordinates = "lon lat" ;
		range_ku:comment = "All instrumental corrections included, i.e. distance antenna-COG (cog_corr), USO drift correction (uso_corr), internal path correction (internal_path_delay_corr_ku), Doppler correction (doppler_corr_ku), modeled instrumental errors correction (modeled_instr_corr_range_ku) and system bias. range updated to account for reference plane and internal path delay " ;
	int range_20hz_ku(time, meas_ind) ;
		range_20hz_ku:_FillValue = 2147483647 ;
		range_20hz_ku:long_name = "20 Hz Ku band corrected altimeter range" ;
		range_20hz_ku:standard_name = "altimeter_range" ;
		range_20hz_ku:units = "m" ;
		range_20hz_ku:add_offset = 1300000. ;
		range_20hz_ku:scale_factor = 0.0001 ;
		range_20hz_ku:coordinates = "lon_20hz lat_20hz" ;
		range_20hz_ku:comment = "All instrumental corrections included, i.e. distance antenna-COG (cog_corr), USO drift correction (uso_corr), internal path correction (internal_path_delay_corr_ku), Doppler correction (doppler_corr_ku), modeled instrumental errors correction (modeled_instr_corr_range_ku) and system bias. range_20hz updated to account for reference plane and internal path delay " ;
	int range_c(time) ;
		range_c:_FillValue = 2147483647 ;
		range_c:long_name = "1 Hz C band corrected altimeter range" ;
		range_c:standard_name = "altimeter_range" ;
		range_c:units = "m" ;
		range_c:quality_flag = "qual_alt_1hz_range_c" ;
		range_c:add_offset = 1300000. ;
		range_c:scale_factor = 0.0001 ;
		range_c:coordinates = "lon lat" ;
		range_c:comment = "All instrumental corrections included, i.e. distance antenna-COG (cog_corr), USO drift correction (uso_corr), internal path correction (internal_path_delay_corr_c), Doppler correction (doppler_corr_c), modeled instrumental errors correction (modeled_instr_corr_range_c) and system bias. range_c updated to account for reference plane and internal path delay " ;
	int range_20hz_c(time, meas_ind) ;
		range_20hz_c:_FillValue = 2147483647 ;
		range_20hz_c:long_name = "20 Hz C band corrected altimeter range" ;
		range_20hz_c:standard_name = "altimeter_range" ;
		range_20hz_c:units = "m" ;
		range_20hz_c:add_offset = 1300000. ;
		range_20hz_c:scale_factor = 0.0001 ;
		range_20hz_c:coordinates = "lon_20hz lat_20hz" ;
		range_20hz_c:comment = "All instrumental corrections included, i.e. distance antenna-COG (cog_corr), USO drift correction (uso_corr), internal path correction (internal_path_delay_corr_c), Doppler correction (doppler_corr_c), modeled instrumental errors correction (modeled_instr_corr_range_c) and system bias. range_20hz_c updated to account for reference plane and internal path delay " ;
	short range_used_20hz_ku(time, meas_ind) ;
		range_used_20hz_ku:_FillValue = 127b ;
		range_used_20hz_ku:long_name = "20 Hz flag for utilization in the computation of 1Hz Ku band range" ;
		range_used_20hz_ku:flag_values = 0b, 1b ;
		range_used_20hz_ku:flag_meanings = "yes no" ;
		range_used_20hz_ku:coordinates = "lon_20hz lat_20hz" ;
		range_used_20hz_ku:comment = "Map of valid points used to compute the 1-Hz Ku-band altimeter range" ;
	short range_used_20hz_c(time, meas_ind) ;
		range_used_20hz_c:_FillValue = 127b ;
		range_used_20hz_c:long_name = "20 Hz flag for utilization in the computation of 1Hz C band range" ;
		range_used_20hz_c:flag_values = 0b, 1b ;
		range_used_20hz_c:flag_meanings = "yes no" ;
		range_used_20hz_c:coordinates = "lon_20hz lat_20hz" ;
		range_used_20hz_c:comment = "Map of valid points used to compute the 1-Hz C-band altimeter range" ;
	short range_rms_ku(time) ;
		range_rms_ku:_FillValue = 32767s ;
		range_rms_ku:long_name = "RMS of the Ku band range" ;
		range_rms_ku:units = "m" ;
		range_rms_ku:scale_factor = 0.0001 ;
		range_rms_ku:coordinates = "lon lat" ;
		range_rms_ku:comment = "Compression of Ku-band high rate elements is preceded by a detection of outliers. Only valid high-rate values are used to compute this element" ;
	short range_rms_c(time) ;
		range_rms_c:_FillValue = 32767s ;
		range_rms_c:long_name = "RMS of the C band range" ;
		range_rms_c:units = "m" ;
		range_rms_c:scale_factor = 0.0001 ;
		range_rms_c:coordinates = "lon lat" ;
		range_rms_c:comment = "Compression of C-band high rate elements is preceded by a detection of outliers. Only valid high-rate values are used to compute this element" ;
	byte range_numval_ku(time) ;
		range_numval_ku:_FillValue = 127b ;
		range_numval_ku:long_name = "number of valid points for Ku band range" ;
		range_numval_ku:units = "count" ;
		range_numval_ku:valid_min = 0b ;
		range_numval_ku:valid_max = 20b ;
		range_numval_ku:coordinates = "lon lat" ;
	byte range_numval_c(time) ;
		range_numval_c:_FillValue = 127b ;
		range_numval_c:long_name = "number of valid points for C band range" ;
		range_numval_c:units = "count" ;
		range_numval_c:valid_min = 0b ;
		range_numval_c:valid_max = 20b ;
		range_numval_c:coordinates = "lon lat" ;
	byte number_of_iterations_ku(time, meas_ind) ;
		number_of_iterations_ku:_FillValue = 127b ;
		number_of_iterations_ku:long_name = "20 Hz number of iterations of the ocean retracking in Ku band" ;
		number_of_iterations_ku:units = "count" ;
		number_of_iterations_ku:coordinates = "lon_20hz lat_20hz" ;
	byte number_of_iterations_c(time, meas_ind) ;
		number_of_iterations_c:_FillValue = 127b ;
		number_of_iterations_c:long_name = "20 Hz number of iterations of the ocean retracking in C band" ;
		number_of_iterations_c:units = "count" ;
		number_of_iterations_c:coordinates = "lon_20hz lat_20hz" ;
	int net_instr_corr_range_ku(time) ;
		net_instr_corr_range_ku:_FillValue = 2147483647 ;
		net_instr_corr_range_ku:long_name = "net instrumental correction on the Ku band range" ;
		net_instr_corr_range_ku:units = "m" ;
		net_instr_corr_range_ku:quality_flag = "qual_inst_corr_1hz_range_ku" ;
		net_instr_corr_range_ku:scale_factor = 0.0001 ;
		net_instr_corr_range_ku:coordinates = "lon lat" ;
		net_instr_corr_range_ku:comment = "Sum of distance antenna-COG (cog_corr), USO drift correction (uso_corr), internal path correction (internal_path_delay_corr_ku), Doppler correction (doppler_corr_ku), modeled instrumental errors correction (modeled_instr_corr_range_ku) and system bias. Updated to account for reference plane and internal path delay " ;
	int net_instr_corr_range_c(time) ;
		net_instr_corr_range_c:_FillValue = 2147483647 ;
		net_instr_corr_range_c:long_name = "net instrumental correction on the C band range" ;
		net_instr_corr_range_c:units = "m" ;
		net_instr_corr_range_c:quality_flag = "qual_inst_corr_1hz_range_c" ;
		net_instr_corr_range_c:scale_factor = 0.0001 ;
		net_instr_corr_range_c:coordinates = "lon lat" ;
		net_instr_corr_range_c:comment = "Sum of distance antenna-COG (cog_corr), USO drift correction (uso_corr), internal path correction (internal_path_delay_corr_c), Doppler correction (doppler_corr_c), modeled instrumental errors correction (modeled_instr_corr_range_c) and system bias. Updated to account for reference plane and internal path delay " ;
	short model_dry_tropo_corr(time) ;
		model_dry_tropo_corr:_FillValue = 32767s ;
		model_dry_tropo_corr:long_name = "model dry tropospheric correction" ;
		model_dry_tropo_corr:standard_name = "altimeter_range_correction_due_to_dry_troposphere" ;
		model_dry_tropo_corr:source = "European Center for Medium Range Weather Forecasting" ;
		model_dry_tropo_corr:institution = "ECMWF" ;
		model_dry_tropo_corr:units = "m" ;
		model_dry_tropo_corr:quality_flag = "" ;
		model_dry_tropo_corr:scale_factor = 0.0001 ;
		model_dry_tropo_corr:coordinates = "lon lat" ;
		model_dry_tropo_corr:comment = "Computed at the altimeter time-tag from the interpolation of 2 meteorological fields that surround the altimeter time-tag. A dry tropospheric correction must be added (negative value) to the instrument range to correct this range measurement for dry tropospheric range delays of the radar pulse. See Jason-1 User Handbook" ;
	short model_dry_tropo_corr_era(time) ;
		model_dry_tropo_corr_era:_FillValue = 32767s ;
		model_dry_tropo_corr_era:long_name = "model dry tropospheric correction from ERA_Interim products" ;
		model_dry_tropo_corr_era:standard_name = "altimeter_range_correction_due_to_dry_troposphere" ;
		model_dry_tropo_corr_era:source = "European Center for Medium Range Weather Forecasting" ;
		model_dry_tropo_corr_era:institution = "ECMWF" ;
		model_dry_tropo_corr_era:units = "m" ;
		model_dry_tropo_corr_era:scale_factor = 0.0001 ;
		model_dry_tropo_corr_era:coordinates = "lon lat" ;
		model_dry_tropo_corr_era:comment = "Courtesy of ECMWF as provider of met data for the atmospheric corrections. Computed at the altimeter time-tag from the interpolation of 2 ERA meteorological fields that surround the altimeter time-tag. A dry tropospheric correction must be added (negative value) to the instrument range to correct this range measurement for dry tropospheric range delays of the radar pulse. See Jason-1 User Handbook" ;
	short model_wet_tropo_corr(time) ;
		model_wet_tropo_corr:_FillValue = 32767s ;
		model_wet_tropo_corr:long_name = "model wet tropospheric correction" ;
		model_wet_tropo_corr:standard_name = "altimeter_range_correction_due_to_wet_troposphere" ;
		model_wet_tropo_corr:source = "European Center for Medium Range Weather Forecasting" ;
		model_wet_tropo_corr:institution = "ECMWF" ;
		model_wet_tropo_corr:units = "m" ;
		model_wet_tropo_corr:quality_flag = "" ;
		model_wet_tropo_corr:scale_factor = 0.0001 ;
		model_wet_tropo_corr:coordinates = "lon lat" ;
		model_wet_tropo_corr:comment = "Computed at the altimeter time-tag from the interpolation of 2 meteorological fields that surround the altimeter time-tag. A wet tropospheric correction must be added (negative value) to the instrument range to correct this range measurement for wet tropospheric range delays of the radar pulse. See Jason-1 User Handbook" ;
	short model_wet_tropo_corr_era(time) ;
		model_wet_tropo_corr_era:_FillValue = 32767s ;
		model_wet_tropo_corr_era:long_name = "model wet tropospheric correction from ERA_Interim products" ;
		model_wet_tropo_corr_era:standard_name = "altimeter_range_correction_due_to_wet_troposphere" ;
		model_wet_tropo_corr_era:source = "European Center for Medium Range Weather Forecasting" ;
		model_wet_tropo_corr_era:institution = "ECMWF" ;
		model_wet_tropo_corr_era:units = "m" ;
		model_wet_tropo_corr_era:scale_factor = 0.0001 ;
		model_wet_tropo_corr_era:coordinates = "lon lat" ;
		model_wet_tropo_corr_era:comment = "Courtesy of ECMWF as provider of met data for the atmospheric corrections. Computed at the altimeter time-tag from the interpolation of 2 ERA meteorological fields that surround the altimeter time-tag. A wet tropospheric correction must be added (negative value) to the instrument range to correct this range measurement for wet tropospheric range delays of the radar pulse. See Jason-1 User Handbook" ;
	short rad_wet_tropo_corr(time) ;
		rad_wet_tropo_corr:_FillValue = 32767s ;
		rad_wet_tropo_corr:long_name = "radiometer wet tropospheric correction" ;
		rad_wet_tropo_corr:standard_name = "altimeter_range_correction_due_to_wet_troposphere" ;
		rad_wet_tropo_corr:source = "JMR" ;
		rad_wet_tropo_corr:institution = "NASA/JPL" ;
		rad_wet_tropo_corr:units = "m" ;
		rad_wet_tropo_corr:quality_flag = "qual_rad_1hz_tb187 and qual_rad_1hz_tb238 and qual_rad_1hz_tb340 and interp_flag_tb" ;
		rad_wet_tropo_corr:scale_factor = 0.0001 ;
		rad_wet_tropo_corr:coordinates = "lon lat" ;
		rad_wet_tropo_corr:comment = "A wet tropospheric correction must be added (negative value) to the instrument range to correct this range measurement for wet tropospheric range delays of the radar pulse" ;
	short iono_corr_alt_ku(time) ;
		iono_corr_alt_ku:_FillValue = 32767s ;
		iono_corr_alt_ku:long_name = "altimeter ionospheric correction on Ku band" ;
		iono_corr_alt_ku:standard_name = "altimeter_range_correction_due_to_ionosphere" ;
		iono_corr_alt_ku:source = "Poseidon-2" ;
		iono_corr_alt_ku:institution = "CNES" ;
		iono_corr_alt_ku:units = "m" ;
		iono_corr_alt_ku:scale_factor = 0.0001 ;
		iono_corr_alt_ku:coordinates = "lon lat" ;
		iono_corr_alt_ku:comment = "An ionospheric correction must be added (negative value) to the instrument range to correct this range measurement for ionospheric range delays of the radar pulse. See Jason-1 User Handbook" ;
	short iono_corr_gim_ku(time) ;
		iono_corr_gim_ku:_FillValue = 32767s ;
		iono_corr_gim_ku:long_name = "GIM ionospheric correction on Ku band" ;
		iono_corr_gim_ku:standard_name = "altimeter_range_correction_due_to_ionosphere" ;
		iono_corr_gim_ku:institution = "NASA/JPL" ;
		iono_corr_gim_ku:units = "m" ;
		iono_corr_gim_ku:scale_factor = 0.0001 ;
		iono_corr_gim_ku:coordinates = "lon lat" ;
		iono_corr_gim_ku:comment = "An ionospheric correction must be added (negative value) to the instrument range to correct this range measurement for ionospheric range delays of the radar pulse. See Jason-1 User Handbook" ;
	short sea_state_bias_ku(time) ;
		sea_state_bias_ku:_FillValue = 32767s ;
		sea_state_bias_ku:long_name = "sea state bias correction in Ku band" ;
		sea_state_bias_ku:standard_name = "sea_surface_height_bias_due_to_sea_surface_roughness" ;
		sea_state_bias_ku:source = "Empirical solution fitted to Jason-1 GDR-C data. Computed using updated values of sigma0 (atmospheric correction being updated)" ;
		sea_state_bias_ku:institution = "CNES" ;
		sea_state_bias_ku:units = "m" ;
		sea_state_bias_ku:scale_factor = 0.0001 ;
		sea_state_bias_ku:coordinates = "lon lat" ;
		sea_state_bias_ku:comment = "Computed using wind speed from sigma0 using updated atmospheric attenuation values. A sea state bias correction must be added (negative value) to the instrument range to correct this range measurement for sea state delays of the radar pulse. This element should not be used over land. See Jason-1 User Handbook" ;
	short sea_state_bias_c(time) ;
		sea_state_bias_c:_FillValue = 32767s ;
		sea_state_bias_c:long_name = "sea state bias correction in C band" ;
		sea_state_bias_c:standard_name = "sea_surface_height_bias_due_to_sea_surface_roughness" ;
		sea_state_bias_c:source = "Empirical solution fitted to Jason-1 GDR-C data. Computed using updated values of sigma0 (atmospheric correction being updated)" ;
		sea_state_bias_c:institution = "CNES" ;
		sea_state_bias_c:units = "m" ;
		sea_state_bias_c:scale_factor = 0.0001 ;
		sea_state_bias_c:coordinates = "lon lat" ;
		sea_state_bias_c:comment = "Computed using wind speed from sigma0 using updated atmospheric attenuation values. A sea state bias correction must be added (negative value) to the instrument range to correct this range measurement for sea state delays of the radar pulse. This element should not be used over land. See Jason-1 User Handbook" ;
	short swh_ku(time) ;
		swh_ku:_FillValue = 32767s ;
		swh_ku:long_name = "Ku band corrected significant waveheight" ;
		swh_ku:standard_name = "sea_surface_wave_significant_height" ;
		swh_ku:units = "m" ;
		swh_ku:quality_flag = "qual_alt_1hz_swh_ku" ;
		swh_ku:scale_factor = 0.001 ;
		swh_ku:coordinates = "lon lat" ;
		swh_ku:comment = "All instrumental corrections included, i.e. modeled instrumental errors correction (modeled_instr_corr_swh_ku) and system bias" ;
	short swh_20hz_ku(time, meas_ind) ;
		swh_20hz_ku:_FillValue = 32767s ;
		swh_20hz_ku:long_name = "20 Hz Ku band corrected significant waveheight" ;
		swh_20hz_ku:standard_name = "sea_surface_wave_significant_height" ;
		swh_20hz_ku:units = "m" ;
		swh_20hz_ku:scale_factor = 0.001 ;
		swh_20hz_ku:coordinates = "lon_20hz lat_20hz" ;
		swh_20hz_ku:comment = "All instrumental corrections included, i.e. modeled instrumental errors correction (modeled_instr_corr_swh_ku) and system bias" ;
	short swh_c(time) ;
		swh_c:_FillValue = 32767s ;
		swh_c:long_name = "C band corrected significant waveheight" ;
		swh_c:standard_name = "sea_surface_wave_significant_height" ;
		swh_c:units = "m" ;
		swh_c:quality_flag = "qual_alt_1hz_swh_c" ;
		swh_c:scale_factor = 0.001 ;
		swh_c:coordinates = "lon lat" ;
		swh_c:comment = "All instrumental corrections included, i.e. modeled instrumental errors correction (modeled_instr_corr_swh_c) and system bias" ;
	short swh_20hz_c(time, meas_ind) ;
		swh_20hz_c:_FillValue = 32767s ;
		swh_20hz_c:long_name = "20 Hz C band corrected significant waveheight" ;
		swh_20hz_c:standard_name = "sea_surface_wave_significant_height" ;
		swh_20hz_c:units = "m" ;
		swh_20hz_c:scale_factor = 0.001 ;
		swh_20hz_c:coordinates = "lon_20hz lat_20hz" ;
		swh_20hz_c:comment = "All instrumental corrections included, i.e. modeled instrumental errors correction (modeled_instr_corr_swh_c) and system bias" ;
	short swh_used_20hz_ku(time, meas_ind) ;
		swh_used_20hz_ku:_FillValue = 127b ;
		swh_used_20hz_ku:long_name = "20 Hz flag for utilization in the computation of 1Hz Ku band significant waveheight" ;
		swh_used_20hz_ku:flag_values = 0b, 1b ;
		swh_used_20hz_ku:flag_meanings = "yes no" ;
		swh_used_20hz_ku:coordinates = "lon_20hz lat_20hz" ;
		swh_used_20hz_ku:comment = "Map of valid points used to compute the 1-Hz Ku-band significant waveheight" ;
	short swh_used_20hz_c(time, meas_ind) ;
		swh_used_20hz_c:_FillValue = 127b ;
		swh_used_20hz_c:long_name = "20 Hz flag for utilization in the computation of 1Hz C band significant waveheight" ;
		swh_used_20hz_c:flag_values = 0b, 1b ;
		swh_used_20hz_c:flag_meanings = "yes no" ;
		swh_used_20hz_c:coordinates = "lon_20hz lat_20hz" ;
		swh_used_20hz_c:comment = "Map of valid points used to compute the 1-Hz C-band significant waveheight" ;
	short swh_rms_ku(time) ;
		swh_rms_ku:_FillValue = 32767s ;
		swh_rms_ku:long_name = "RMS of the Ku band significant waveheight" ;
		swh_rms_ku:units = "m" ;
		swh_rms_ku:scale_factor = 0.001 ;
		swh_rms_ku:coordinates = "lon lat" ;
		swh_rms_ku:comment = "Compression of Ku-band high rate elements is preceded by a detection of outliers. Only valid high-rate values are used to compute this element" ;
	short swh_rms_c(time) ;
		swh_rms_c:_FillValue = 32767s ;
		swh_rms_c:long_name = "RMS of the C band significant waveheight" ;
		swh_rms_c:units = "m" ;
		swh_rms_c:scale_factor = 0.001 ;
		swh_rms_c:coordinates = "lon lat" ;
		swh_rms_c:comment = "Compression of C-band high rate elements is preceded by a detection of outliers. Only valid high-rate values are used to compute this element" ;
	short swh_numval_ku(time) ;
		swh_numval_ku:_FillValue = 127b ;
		swh_numval_ku:long_name = "number of valid points used to compute Ku significant waveheight" ;
		swh_numval_ku:units = "count" ;
		swh_numval_ku:valid_min = 0b ;
		swh_numval_ku:valid_max = 20b ;
		swh_numval_ku:coordinates = "lon lat" ;
	short swh_numval_c(time) ;
		swh_numval_c:_FillValue = 127b ;
		swh_numval_c:long_name = "number of valid points used to compute C significant waveheight" ;
		swh_numval_c:units = "count" ;
		swh_numval_c:valid_min = 0b ;
		swh_numval_c:valid_max = 20b ;
		swh_numval_c:coordinates = "lon lat" ;
	short net_instr_corr_swh_ku(time) ;
		net_instr_corr_swh_ku:_FillValue = 32767s ;
		net_instr_corr_swh_ku:long_name = "net instrumental correction on Ku band significant waveheight" ;
		net_instr_corr_swh_ku:units = "m" ;
		net_instr_corr_swh_ku:quality_flag = "qual_inst_corr_1hz_swh_ku" ;
		net_instr_corr_swh_ku:scale_factor = 0.001 ;
		net_instr_corr_swh_ku:coordinates = "lon lat" ;
		net_instr_corr_swh_ku:comment = "Sum of modeled instrumental errors correction (modeled_instr_corr_swh_ku) and system bias" ;
	short net_instr_corr_swh_c(time) ;
		net_instr_corr_swh_c:_FillValue = 32767s ;
		net_instr_corr_swh_c:long_name = "net instrumental correction on C band significant waveheight" ;
		net_instr_corr_swh_c:units = "m" ;
		net_instr_corr_swh_c:quality_flag = "qual_inst_corr_1hz_swh_c" ;
		net_instr_corr_swh_c:scale_factor = 0.001 ;
		net_instr_corr_swh_c:coordinates = "lon lat" ;
		net_instr_corr_swh_c:comment = "Sum of modeled instrumental errors correction (modeled_instr_corr_swh_c) and system bias" ;
	short sig0_ku(time) ;
		sig0_ku:_FillValue = 32767s ;
		sig0_ku:long_name = "Ku band corrected backscatter coefficient" ;
		sig0_ku:standard_name = "surface_backwards_scattering_coefficient_of_radar_wave" ;
		sig0_ku:units = "dB" ;
		sig0_ku:quality_flag = "qual_alt_1hz_sig0_ku" ;
		sig0_ku:scale_factor = 0.01 ;
		sig0_ku:coordinates = "lon lat" ;
		sig0_ku:comment = "All instrumental corrections included, excepted the system bias, i.e. AGC instrumental errors correction, internal calibration correction (internal_corr_sig0_ku), modeled instrumental errors correction (modeled_instr_corr_sig0_ku) and atmospheric attenuation (atmos_corr_sig0_ku)" ;
	short sig0_20hz_ku(time, meas_ind) ;
		sig0_20hz_ku:_FillValue = 32767s ;
		sig0_20hz_ku:long_name = "20 Hz Ku band corrected backscatter coefficient" ;
		sig0_20hz_ku:standard_name = "surface_backwards_scattering_coefficient_of_radar_wave" ;
		sig0_20hz_ku:units = "dB" ;
		sig0_20hz_ku:scale_factor = 0.01 ;
		sig0_20hz_ku:coordinates = "lon_20hz lat_20hz" ;
		sig0_20hz_ku:comment = "All instrumental corrections included, excepted the system bias, i.e. AGC instrumental errors correction, internal calibration correction (internal_corr_sig0_ku), modeled instrumental errors correction (modeled_instr_corr_sig0_ku) and atmospheric attenuation (atmos_corr_sig0_ku)" ;
	short sig0_c(time) ;
		sig0_c:_FillValue = 32767s ;
		sig0_c:long_name = "C band corrected backscatter coefficient" ;
		sig0_c:standard_name = "surface_backwards_scattering_coefficient_of_radar_wave" ;
		sig0_c:units = "dB" ;
		sig0_c:quality_flag = "qual_alt_1hz_sig0_c" ;
		sig0_c:scale_factor = 0.01 ;
		sig0_c:coordinates = "lon lat" ;
		sig0_c:comment = "All instrumental corrections included, excepted the system bias, i.e. AGC instrumental errors correction, internal calibration correction (internal_corr_sig0_c), modeled instrumental errors correction (modeled_instr_corr_sig0_c) and atmospheric attenuation (atmos_corr_sig0_c)" ;
	short sig0_20hz_c(time, meas_ind) ;
		sig0_20hz_c:_FillValue = 32767s ;
		sig0_20hz_c:long_name = "20 Hz C band corrected backscatter coefficient" ;
		sig0_20hz_c:standard_name = "surface_backwards_scattering_coefficient_of_radar_wave" ;
		sig0_20hz_c:units = "dB" ;
		sig0_20hz_c:scale_factor = 0.01 ;
		sig0_20hz_c:coordinates = "lon_20hz lat_20hz" ;
		sig0_20hz_c:comment = "All instrumental corrections included, excepted the system bias, i.e. AGC instrumental errors correction, internal calibration correction (internal_corr_sig0_c), modeled instrumental errors correction (modeled_instr_corr_sig0_c) and atmospheric attenuation (atmos_corr_sig0_c)" ;
	byte sig0_used_20hz_ku(time, meas_ind) ;
		sig0_used_20hz_ku:_FillValue = 127b ;
		sig0_used_20hz_ku:long_name = "20 Hz flag for utilization in the computation of 1Hz Ku band backscatter coefficient" ;
		sig0_used_20hz_ku:flag_values = 0b, 1b ;
		sig0_used_20hz_ku:flag_meanings = "yes no" ;
		sig0_used_20hz_ku:coordinates = "lon_20hz lat_20hz" ;
		sig0_used_20hz_ku:comment = "Map of valid points used to compute the 1-Hz Ku-band backscatter coefficient" ;
	byte sig0_used_20hz_c(time, meas_ind) ;
		sig0_used_20hz_c:_FillValue = 127b ;
		sig0_used_20hz_c:long_name = "20 Hz flag for utilization in the computation of 1Hz C band backscatter coefficient" ;
		sig0_used_20hz_c:flag_values = 0b, 1b ;
		sig0_used_20hz_c:flag_meanings = "yes no" ;
		sig0_used_20hz_c:coordinates = "lon_20hz lat_20hz" ;
		sig0_used_20hz_c:comment = "Map of valid points used to compute the 1-Hz C-band backscatter coefficient" ;
	short sig0_rms_ku(time) ;
		sig0_rms_ku:_FillValue = 32767s ;
		sig0_rms_ku:long_name = "RMS of the Ku band backscatter coefficient" ;
		sig0_rms_ku:units = "dB" ;
		sig0_rms_ku:scale_factor = 0.01 ;
		sig0_rms_ku:coordinates = "lon lat" ;
		sig0_rms_ku:comment = "Compression of Ku-band high rate elements is preceded by a detection of outliers. Only valid high-rate values are used to compute this element" ;
	short sig0_rms_c(time) ;
		sig0_rms_c:_FillValue = 32767s ;
		sig0_rms_c:long_name = "RMS of the C band backscatter coefficient" ;
		sig0_rms_c:units = "dB" ;
		sig0_rms_c:scale_factor = 0.01 ;
		sig0_rms_c:coordinates = "lon lat" ;
		sig0_rms_c:comment = "Compression of C-band high rate elements is preceded by a detection of outliers. Only valid high-rate values are used to compute this element" ;
	byte sig0_numval_ku(time) ;
		sig0_numval_ku:_FillValue = 127b ;
		sig0_numval_ku:long_name = "number of valid points used to compute Ku backscatter coefficient" ;
		sig0_numval_ku:units = "count" ;
		sig0_numval_ku:valid_min = 0b ;
		sig0_numval_ku:valid_max = 20b ;
		sig0_numval_ku:coordinates = "lon lat" ;
	byte sig0_numval_c(time) ;
		sig0_numval_c:_FillValue = 127b ;
		sig0_numval_c:long_name = "number of valid points used to compute C backscatter coefficient" ;
		sig0_numval_c:units = "count" ;
		sig0_numval_c:valid_min = 0b ;
		sig0_numval_c:valid_max = 20b ;
		sig0_numval_c:coordinates = "lon lat" ;
	short agc_ku(time) ;
		agc_ku:_FillValue = 32767s ;
		agc_ku:long_name = "Ku band corrected AGC" ;
		agc_ku:units = "dB" ;
		agc_ku:scale_factor = 0.01 ;
		agc_ku:coordinates = "lon lat" ;
		agc_ku:comment = "AGC is corrected for instrumental errors due to the imperfections of the on-board attenuators" ;
	short agc_c(time) ;
		agc_c:_FillValue = 32767s ;
		agc_c:long_name = "C band corrected AGC" ;
		agc_c:units = "dB" ;
		agc_c:scale_factor = 0.01 ;
		agc_c:coordinates = "lon lat" ;
		agc_c:comment = "AGC is corrected for instrumental errors due to the imperfections of the on-board attenuators" ;
	short agc_rms_ku(time) ;
		agc_rms_ku:_FillValue = 32767s ;
		agc_rms_ku:long_name = "RMS of the Ku band AGC" ;
		agc_rms_ku:units = "dB" ;
		agc_rms_ku:scale_factor = 0.01 ;
		agc_rms_ku:coordinates = "lon lat" ;
		agc_rms_ku:comment = "Compression of Ku-band high rate elements is preceded by a detection of outliers. Only valid high-rate values are used to compute this element" ;
	short agc_rms_c(time) ;
		agc_rms_c:_FillValue = 32767s ;
		agc_rms_c:long_name = "RMS of the C band AGC" ;
		agc_rms_c:units = "dB" ;
		agc_rms_c:scale_factor = 0.01 ;
		agc_rms_c:coordinates = "lon lat" ;
		agc_rms_c:comment = "Compression of C-band high rate elements is preceded by a detection of outliers. Only valid high-rate values are used to compute this element" ;
	byte agc_numval_ku(time) ;
		agc_numval_ku:_FillValue = 127b ;
		agc_numval_ku:long_name = "number of valid points used to compute Ku band AGC" ;
		agc_numval_ku:units = "count" ;
		agc_numval_ku:valid_min = 0b ;
		agc_numval_ku:valid_max = 20b ;
		agc_numval_ku:coordinates = "lon lat" ;
	byte agc_numval_c(time) ;
		agc_numval_c:_FillValue = 127b ;
		agc_numval_c:long_name = "number of valid points used to compute C band AGC" ;
		agc_numval_c:units = "count" ;
		agc_numval_c:valid_min = 0b ;
		agc_numval_c:valid_max = 20b ;
		agc_numval_c:coordinates = "lon lat" ;
	short net_instr_corr_sig0_ku(time) ;
		net_instr_corr_sig0_ku:_FillValue = 32767s ;
		net_instr_corr_sig0_ku:long_name = "net instrumental correction on Ku backscatter coefficient" ;
		net_instr_corr_sig0_ku:units = "dB" ;
		net_instr_corr_sig0_ku:quality_flag = "qual_inst_corr_1hz_sig0_ku" ;
		net_instr_corr_sig0_ku:scale_factor = 0.01 ;
		net_instr_corr_sig0_ku:coordinates = "lon lat" ;
		net_instr_corr_sig0_ku:comment = "Sum of AGC instrumental errors correction, internal calibration correction (internal_corr_sig0_ku) and modeled instrumental errors correction (modeled_instr_corr_sig0_ku) - system bias not included" ;
	short net_instr_corr_sig0_c(time) ;
		net_instr_corr_sig0_c:_FillValue = 32767s ;
		net_instr_corr_sig0_c:long_name = "net instrumental correction on C backscatter coefficient" ;
		net_instr_corr_sig0_c:units = "dB" ;
		net_instr_corr_sig0_c:quality_flag = "qual_inst_corr_1hz_sig0_c" ;
		net_instr_corr_sig0_c:scale_factor = 0.01 ;
		net_instr_corr_sig0_c:coordinates = "lon lat" ;
		net_instr_corr_sig0_c:comment = "Sum of AGC instrumental errors correction, internal calibration correction (internal_corr_sig0_c) and modeled instrumental errors correction (modeled_instr_corr_sig0_c) - system bias not included" ;
	short atmos_corr_sig0_ku(time) ;
		atmos_corr_sig0_ku:_FillValue = 32767s ;
		atmos_corr_sig0_ku:long_name = "atmospheric attenuation correction on Ku band backscatter coefficient" ;
		atmos_corr_sig0_ku:units = "dB" ;
		atmos_corr_sig0_ku:scale_factor = 0.01 ;
		atmos_corr_sig0_ku:coordinates = "lon lat" ;
	short atmos_corr_sig0_c(time) ;
		atmos_corr_sig0_c:_FillValue = 32767s ;
		atmos_corr_sig0_c:long_name = "atmospheric attenuation correction on C band backscatter coefficient" ;
		atmos_corr_sig0_c:units = "dB" ;
		atmos_corr_sig0_c:scale_factor = 0.01 ;
		atmos_corr_sig0_c:coordinates = "lon lat" ;
	short off_nadir_angle_wf_ku(time) ;
		off_nadir_angle_wf_ku:_FillValue = 32767s ;
		off_nadir_angle_wf_ku:long_name = "square of the off nadir angle computed from Ku waveforms" ;
		off_nadir_angle_wf_ku:units = "degrees^2" ;
		off_nadir_angle_wf_ku:quality_flag = "qual_alt_1hz_off_nadir_angle_wf_ku" ;
		off_nadir_angle_wf_ku:scale_factor = 0.0001 ;
		off_nadir_angle_wf_ku:coordinates = "lon lat" ;
	short tb_187(time) ;
		tb_187:_FillValue = 32767s ;
		tb_187:long_name = "18.7 GHz main beam brightness temperature" ;
		tb_187:standard_name = "surface_brightness_temperature" ;
		tb_187:units = "K" ;
		tb_187:quality_flag = "qual_rad_1hz_tb187" ;
		tb_187:scale_factor = 0.01 ;
		tb_187:coordinates = "lon lat" ;
		tb_187:comment = "Brightness temperatures are unsmoothed (along-track averaging has not been performed on the brightness temperatures)" ;
	short tb_238(time) ;
		tb_238:_FillValue = 32767s ;
		tb_238:long_name = "23.8 GHz main beam brightness temperature" ;
		tb_238:standard_name = "surface_brightness_temperature" ;
		tb_238:units = "K" ;
		tb_238:quality_flag = "qual_rad_1hz_tb238" ;
		tb_238:scale_factor = 0.01 ;
		tb_238:coordinates = "lon lat" ;
		tb_238:comment = "Brightness temperatures are unsmoothed (along-track averaging has not been performed on the brightness temperatures)" ;
	short tb_340(time) ;
		tb_340:_FillValue = 32767s ;
		tb_340:long_name = "34.0 GHz main beam brightness temperature" ;
		tb_340:standard_name = "surface_brightness_temperature" ;
		tb_340:units = "K" ;
		tb_340:quality_flag = "qual_rad_1hz_tb340" ;
		tb_340:scale_factor = 0.01 ;
		tb_340:coordinates = "lon lat" ;
		tb_340:comment = "Brightness temperatures are unsmoothed (along-track averaging has not been performed on the brightness temperatures)" ;
	short tb_187_smoothed(time) ;
		tb_187_smoothed:_FillValue = 32767s ;
		tb_187_smoothed:long_name = "18.7 GHz main beam smoothed brightness temperature" ;
		tb_187_smoothed:standard_name = "surface_brightness_temperature" ;
		tb_187_smoothed:units = "K" ;
		tb_187_smoothed:quality_flag = "qual_rad_1hz_tb187" ;
		tb_187_smoothed:scale_factor = 0.01 ;
		tb_187_smoothed:coordinates = "lon lat" ;
		tb_187_smoothed:comment = "Brightness temperatures are along-track averaged" ;
	short tb_238_smoothed(time) ;
		tb_238_smoothed:_FillValue = 32767s ;
		tb_238_smoothed:long_name = "23.8 GHz main beam smoothed brightness temperature" ;
		tb_238_smoothed:standard_name = "surface_brightness_temperature" ;
		tb_238_smoothed:units = "K" ;
		tb_238_smoothed:quality_flag = "qual_rad_1hz_tb238" ;
		tb_238_smoothed:scale_factor = 0.01 ;
		tb_238_smoothed:coordinates = "lon lat" ;
		tb_238_smoothed:comment = "Brightness temperatures are along-track averaged" ;
	short tb_340_smoothed(time) ;
		tb_340_smoothed:_FillValue = 32767s ;
		tb_340_smoothed:long_name = "34.0 GHz main beam smoothed brightness temperature" ;
		tb_340_smoothed:standard_name = "surface_brightness_temperature" ;
		tb_340_smoothed:units = "K" ;
		tb_340_smoothed:quality_flag = "qual_rad_1hz_tb340" ;
		tb_340_smoothed:scale_factor = 0.01 ;
		tb_340_smoothed:coordinates = "lon lat" ;
		tb_340_smoothed:comment = "Brightness temperatures are along-track averaged" ;
	int mean_sea_surface(time) ;
		mean_sea_surface:_FillValue = 2147483647 ;
		mean_sea_surface:long_name = "mean sea surface height above reference ellipsoid" ;
		mean_sea_surface:source = "MSS_CNES_CLS-2011" ;
		mean_sea_surface:institution = "CLS/CNES" ;
		mean_sea_surface:units = "m" ;
		mean_sea_surface:quality_flag = "mean_sea_surface_err" ;
		mean_sea_surface:scale_factor = 0.0001 ;
		mean_sea_surface:coordinates = "lon lat" ;
		mean_sea_surface:comment = "The mean sea surface height is referenced to a 20 years mean. See Jason-1 User Handbook." ;
	int mean_sea_surface_err(time) ;
		mean_sea_surface_err:_FillValue = 2147483647 ;
		mean_sea_surface_err:long_name = "calibrated error of mean sea surface" ;
		mean_sea_surface_err:source = "MSS_CNES_CLS-2011" ;
		mean_sea_surface_err:institution = "CLS/CNES" ;
		mean_sea_surface_err:units = "m" ;
		mean_sea_surface_err:scale_factor = 0.0001 ;
		mean_sea_surface_err:coordinates = "lon lat" ;
		mean_sea_surface_err:comment = "See Jason-1 User Handbook" ;
	int mean_topography(time) ;
		mean_topography:_FillValue = 2147483647 ;
		mean_topography:long_name = "mean dynamic topography above geoid" ;
		mean_topography:source = "MDT_CNES_CLS-2013" ;
		mean_topography:institution = "CLS/CNES" ;
		mean_topography:units = "m" ;
		mean_topography:quality_flag = "mean_topography_err" ;
		mean_topography:scale_factor = 0.0001 ;
		mean_topography:coordinates = "lon lat" ;
		mean_topography:comment = "The mean dynamic topography is referenced to a 20 years mean. See Jason-1 User Handbook." ;
	int mean_topography_err(time) ;
		mean_topography_err:_FillValue = 2147483647 ;
		mean_topography_err:long_name = "error on mean dynamic topography" ;
		mean_topography_err:source = "MDT_CNES_CLS-2013" ;
		mean_topography_err:institution = "CLS/CNES" ;
		mean_topography_err:units = "m" ;
		mean_topography_err:scale_factor = 0.0001 ;
		mean_topography_err:coordinates = "lon lat" ;
		mean_topography_err:comment = "See Jason-1 User Handbook" ;
	int geoid(time) ;
		geoid:_FillValue = 2147483647 ;
		geoid:long_name = "geoid height" ;
		geoid:standard_name = "geoid_height_above_reference_ellipsoid" ;
		geoid:source = "EGM2008" ;
		geoid:institution = "National Geospatial-Intelligence Agency (NGA)" ;
		geoid:units = "m" ;
		geoid:scale_factor = 0.0001 ;
		geoid:coordinates = "lon lat" ;
		geoid:comment = "Computed from the geoid model with a correction to refer the value to the mean tide system i.e. includes the permanent tide (zero frequency). See Jason-1 User Handbook" ;
	int bathymetry(time) ;
		bathymetry:_FillValue = 2147483647 ;
		bathymetry:long_name = "ocean depth/land elevation" ;
		bathymetry:source = "DTM2000.1" ;
		bathymetry:institution = "GSFC" ;
		bathymetry:units = "m" ;
		bathymetry:coordinates = "lon lat" ;
	short inv_bar_corr(time) ;
		inv_bar_corr:_FillValue = 32767s ;
		inv_bar_corr:long_name = "inverted barometer height correction" ;
		inv_bar_corr:standard_name = "sea_surface_height_correction_due_to_air_pressure_at_low_frequency" ;
		inv_bar_corr:source = "European Center for Medium Range Weather Forecasting" ;
		inv_bar_corr:institution = "ECMWF" ;
		inv_bar_corr:units = "m" ;
		inv_bar_corr:quality_flag = "" ;
		inv_bar_corr:scale_factor = 0.0001 ;
		inv_bar_corr:coordinates = "lon lat" ;
		inv_bar_corr:comment = "Computed at the altimeter time-tag from the interpolation of 2 meteorological fields that surround the altimeter time-tag. See Jason-1 User Handbook" ;
	short hf_fluctuations_corr(time) ;
		hf_fluctuations_corr:_FillValue = 32767s ;
		hf_fluctuations_corr:long_name = "high frequency fluctuations of the sea surface topography" ;
		hf_fluctuations_corr:standard_name = "sea_surface_height_correction_due_to_air_pressure_and_wind_at_high_frequency" ;
		hf_fluctuations_corr:institution = "LEGOS/CLS/CNES" ;
		hf_fluctuations_corr:units = "m" ;
		hf_fluctuations_corr:scale_factor = 0.0001 ;
		hf_fluctuations_corr:coordinates = "lon lat" ;
		hf_fluctuations_corr:comment = "Provided as a correction to the inverted barometer correction (inv_bar_corr)" ;
	short inv_bar_corr_era(time) ;
		inv_bar_corr_era:_FillValue = 32767s ;
		inv_bar_corr_era:long_name = "inverted barometer height correction from ERA_Interim products" ;
		inv_bar_corr_era:standard_name = "sea_surface_height_correction_due_to_air_pressure_at_low_frequency" ;
		inv_bar_corr_era:source = "European Center for Medium Range Weather Forecasting" ;
		inv_bar_corr_era:institution = "ECMWF" ;
		inv_bar_corr_era:units = "m" ;
		inv_bar_corr_era:scale_factor = 0.0001 ;
		inv_bar_corr_era:coordinates = "lon lat" ;
		inv_bar_corr_era:comment = "Courtesy of ECMWF as provider of met data for the atmospheric corrections. Computed at the altimeter time-tag from the interpolation of 2 meteorological fields that surround the altimeter time-tag. See Jason-1 User Handbook" ;
	short hf_fluctuations_corr_era(time) ;
		hf_fluctuations_corr_era:_FillValue = 32767s ;
		hf_fluctuations_corr_era:long_name = "high frequency fluctuations of the sea surface topography derived from ERA_Interim products" ;
		hf_fluctuations_corr_era:standard_name = "sea_surface_height_correction_due_to_air_pressure_and_wind_at_high_frequency" ;
		hf_fluctuations_corr_era:institution = "LEGOS/CLS/CNES" ;
		hf_fluctuations_corr_era:units = "m" ;
		hf_fluctuations_corr_era:scale_factor = 0.0001 ;
		hf_fluctuations_corr_era:coordinates = "lon lat" ;
		hf_fluctuations_corr_era:comment = "Provided as a correction to the inverted barometer correction from ERA_Interim products (inv_bar_corr_era)" ;
	int ocean_tide_sol1(time) ;
		ocean_tide_sol1:_FillValue = 2147483647 ;
		ocean_tide_sol1:long_name = "geocentric ocean tide height (solution 1)" ;
		ocean_tide_sol1:standard_name = "sea_surface_height_amplitude_due_to_geocentric_ocean_tide" ;
		ocean_tide_sol1:source = "GOT4.10" ;
		ocean_tide_sol1:institution = "GSFC" ;
		ocean_tide_sol1:units = "m" ;
		ocean_tide_sol1:quality_flag = "interp_flag_ocean_tide_sol1" ;
		ocean_tide_sol1:scale_factor = 0.0001 ;
		ocean_tide_sol1:coordinates = "lon lat" ;
		ocean_tide_sol1:comment = "Solution 1 corresponds to GOT4.10 model. Includes the corresponding loading tide (load_tide_sol1) and equilibrium long-period ocean tide height (ocean_tide_equil). The permanent tide (zero frequency) is not included in this parameter because it is included in the geoid and mean sea surface (geoid, mean_sea_surface). See Jason-1 User Handbook" ;
	int ocean_tide_sol2(time) ;
		ocean_tide_sol2:_FillValue = 2147483647 ;
		ocean_tide_sol2:long_name = "geocentric ocean tide height (solution 2)" ;
		ocean_tide_sol2:standard_name = "sea_surface_height_amplitude_due_to_geocentric_ocean_tide" ;
		ocean_tide_sol2:source = "FES2014" ;
		ocean_tide_sol2:institution = "LEGOS/CNES" ;
		ocean_tide_sol2:units = "m" ;
		ocean_tide_sol2:quality_flag = "interp_flag_ocean_tide_sol2" ;
		ocean_tide_sol2:scale_factor = 0.0001 ;
		ocean_tide_sol2:coordinates = "lon lat" ;
		ocean_tide_sol2:comment = "Solution 2 corresponds to FES2014 model. Includes the corresponding loading tide (load_tide_sol2) and equilibrium long-period ocean tide height (ocean_tide_equil). The permanent tide (zero frequency) is not included in this parameter because it is included in the geoid and mean sea surface (geoid, mean_sea_surface). See Jason-1 User Handbook" ;
	short ocean_tide_equil(time) ;
		ocean_tide_equil:_FillValue = 32767s ;
		ocean_tide_equil:long_name = "equilibrium long-period ocean tide height" ;
		ocean_tide_equil:standard_name = "sea_surface_height_amplitude_due_to_equilibrium_ocean_tide" ;
		ocean_tide_equil:source = "Cartwright and Edden [1973] Corrected tables of tidal harmonics - J. Geophys. J. R. Astr. Soc., 33, 253-264." ;
		ocean_tide_equil:units = "m" ;
		ocean_tide_equil:scale_factor = 0.0001 ;
		ocean_tide_equil:coordinates = "lon lat" ;
		ocean_tide_equil:comment = "This value has already been added to the two geocentric ocean tide height values recorded in the product (ocean_tide_sol1 and ocean_tide_sol2). The permanent tide (zero frequency) is not included in this parameter because it is included in the geoid and mean sea surface (geoid, mean_sea_surface). See Jason-1 User Handbook" ;
	short ocean_tide_non_equil(time) ;
		ocean_tide_non_equil:_FillValue = 32767s ;
		ocean_tide_non_equil:long_name = "non-equilibrium long-period ocean tide height" ;
		ocean_tide_non_equil:standard_name = "sea_surface_height_amplitude_due_to_non_equilibrium_ocean_tide" ;
		ocean_tide_non_equil:source = "FES2014" ;
		ocean_tide_non_equil:institution = "LEGOS/CNES" ;
		ocean_tide_non_equil:units = "m" ;
		ocean_tide_non_equil:scale_factor = 0.0001 ;
		ocean_tide_non_equil:coordinates = "lon lat" ;
		ocean_tide_non_equil:comment = "This parameter is computed as a correction to the parameter ocean_tide_equil. This value can be added to ocean_tide_equil (or ocean_tide_sol1, ocean_tide_sol2) so that the resulting value models the total non equilibrium ocean tide height. See Jason-1 User Handbook" ;
	short load_tide_sol1(time) ;
		load_tide_sol1:_FillValue = 32767s ;
		load_tide_sol1:long_name = "load tide height for geocentric ocean tide (solution 1)" ;
		load_tide_sol1:source = "GOT4.10" ;
		load_tide_sol1:institution = "GSFC" ;
		load_tide_sol1:units = "m" ;
		load_tide_sol1:scale_factor = 0.0001 ;
		load_tide_sol1:coordinates = "lon lat" ;
		load_tide_sol1:comment = "This value has already been added to the corresponding ocean tide height value recorded in the product (ocean_tide_sol1). See Jason-1 User Handbook" ;
	short load_tide_sol2(time) ;
		load_tide_sol2:_FillValue = 32767s ;
		load_tide_sol2:long_name = "load tide height for geocentric ocean tide (solution 2)" ;
		load_tide_sol2:source = "GOT4.8ac, tidal geocenter adjustement included" ;
		load_tide_sol2:institution = "GSFC" ;
		load_tide_sol2:units = "m" ;
		load_tide_sol2:scale_factor = 0.0001 ;
		load_tide_sol2:coordinates = "lon lat" ;
		load_tide_sol2:comment = "This value has already been added to the corresponding ocean tide height value recorded in the product (ocean_tide_sol2). See Jason-1 User Handbook" ;
	short solid_earth_tide(time) ;
		solid_earth_tide:_FillValue = 32767s ;
		solid_earth_tide:long_name = "solid earth tide height" ;
		solid_earth_tide:standard_name = "sea_surface_height_amplitude_due_to_earth_tide" ;
		solid_earth_tide:source = "Cartwright and Edden [1973] Corrected tables of tidal harmonics - J. Geophys. J. R. Astr. Soc., 33, 253-264." ;
		solid_earth_tide:units = "m" ;
		solid_earth_tide:scale_factor = 0.0001 ;
		solid_earth_tide:coordinates = "lon lat" ;
		solid_earth_tide:comment = "Calculated using Cartwright and Tayler tables and consisting of the second and third degree constituents. The permanent tide (zero frequency) is not included. See Jason-1 User Handbook" ;
	short pole_tide(time) ;
		pole_tide:_FillValue = 32767s ;
		pole_tide:long_name = "geocentric pole tide height" ;
		pole_tide:standard_name = "sea_surface_height_amplitude_due_to_pole_tide" ;
		pole_tide:source = "Wahr [1985] Deformation of the Earth induced by polar motion - J. Geophys. Res. (Solid Earth), 90, 9363-9368." ;
		pole_tide:units = "m" ;
		pole_tide:scale_factor = 0.0001 ;
		pole_tide:coordinates = "lon lat" ;
		pole_tide:comment = "See Jason-1 User Handbook" ;
	short wind_speed_model_u(time) ;
		wind_speed_model_u:_FillValue = 32767s ;
		wind_speed_model_u:long_name = "U component of the model wind vector" ;
		wind_speed_model_u:standard_name = "wind_speed" ;
		wind_speed_model_u:source = "European Center for Medium Range Weather Forecasting" ;
		wind_speed_model_u:institution = "ECMWF" ;
		wind_speed_model_u:units = "m/s" ;
		wind_speed_model_u:quality_flag = "" ;
		wind_speed_model_u:scale_factor = 0.01 ;
		wind_speed_model_u:coordinates = "lon lat" ;
		wind_speed_model_u:comment = "Computed at the altimeter time-tag from the interpolation of 2 meteorological fields that surround the altimeter time-tag. See Jason-1 User Handbook" ;
	short wind_speed_model_v(time) ;
		wind_speed_model_v:_FillValue = 32767s ;
		wind_speed_model_v:long_name = "V component of the model wind vector" ;
		wind_speed_model_v:standard_name = "wind_speed" ;
		wind_speed_model_v:source = "European Center for Medium Range Weather Forecasting" ;
		wind_speed_model_v:institution = "ECMWF" ;
		wind_speed_model_v:units = "m/s" ;
		wind_speed_model_v:quality_flag = "" ;
		wind_speed_model_v:scale_factor = 0.01 ;
		wind_speed_model_v:coordinates = "lon lat" ;
		wind_speed_model_v:comment = "Computed at the altimeter time-tag from the interpolation of 2 meteorological fields that surround the altimeter time-tag. See Jason-1 User Handbook" ;
	short wind_speed_model_u_era(time) ;
		wind_speed_model_u_era:_FillValue = 32767s ;
		wind_speed_model_u_era:long_name = "U component of the model wind vector from ERA_Interim products" ;
		wind_speed_model_u_era:standard_name = "wind_speed" ;
		wind_speed_model_u_era:source = "European Center for Medium Range Weather Forecasting" ;
		wind_speed_model_u_era:institution = "ECMWF" ;
		wind_speed_model_u_era:units = "m/s" ;
		wind_speed_model_u_era:scale_factor = 0.01 ;
		wind_speed_model_u_era:coordinates = "lon lat" ;
		wind_speed_model_u_era:comment = "Courtesy of ECMWF. Computed at the altimeter time-tag from the interpolation of 2 meteorological fields that surround the altimeter time-tag. See Jason-1 User Handbook" ;
	short wind_speed_model_v_era(time) ;
		wind_speed_model_v_era:_FillValue = 32767s ;
		wind_speed_model_v_era:long_name = "V component of the model wind vector from ERA_Interim products" ;
		wind_speed_model_v_era:standard_name = "wind_speed" ;
		wind_speed_model_v_era:source = "European Center for Medium Range Weather Forecasting" ;
		wind_speed_model_v_era:institution = "ECMWF" ;
		wind_speed_model_v_era:units = "m/s" ;
		wind_speed_model_v_era:scale_factor = 0.01 ;
		wind_speed_model_v_era:coordinates = "lon lat" ;
		wind_speed_model_v_era:comment = "Courtesy of ECMWF. Computed at the altimeter time-tag from the interpolation of 2 meteorological fields that surround the altimeter time-tag. See Jason-1 User Handbook" ;
	short wind_speed_alt(time) ;
		wind_speed_alt:_FillValue = 32767s ;
		wind_speed_alt:long_name = "altimeter wind speed" ;
		wind_speed_alt:standard_name = "wind_speed" ;
		wind_speed_alt:units = "m/s" ;
		wind_speed_alt:scale_factor = 0.01 ;
		wind_speed_alt:coordinates = "lon lat" ;
		wind_speed_alt:comment = "Should not be used over land. See Jason-1 User Handbook " ;
	short wind_speed_rad(time) ;
		wind_speed_rad:_FillValue = 32767s ;
		wind_speed_rad:long_name = "radiometer wind speed" ;
		wind_speed_rad:standard_name = "wind_speed" ;
		wind_speed_rad:source = "JMR" ;
		wind_speed_rad:institution = "NASA/JPL" ;
		wind_speed_rad:units = "m/s" ;
		wind_speed_rad:scale_factor = 0.01 ;
		wind_speed_rad:coordinates = "lon lat" ;
		wind_speed_rad:comment = "Should not be used over land. See Jason-1 User Handbook" ;
	short rad_water_vapor(time) ;
		rad_water_vapor:_FillValue = 32767s ;
		rad_water_vapor:long_name = "radiometer water vapor content" ;
		rad_water_vapor:standard_name = "atmosphere_water_vapor_content" ;
		rad_water_vapor:source = "JMR" ;
		rad_water_vapor:institution = "NASA/JPL" ;
		rad_water_vapor:units = "kg/m^2" ;
		rad_water_vapor:quality_flag = "qual_rad_1hz_tb187 and qual_rad_1hz_tb238 and qual_rad_1hz_tb340 and interp_flag_tb" ;
		rad_water_vapor:scale_factor = 0.1 ;
		rad_water_vapor:coordinates = "lon lat" ;
		rad_water_vapor:comment = "Should not be used over land." ;
	short rad_liquid_water(time) ;
		rad_liquid_water:_FillValue = 32767s ;
		rad_liquid_water:long_name = "radiometer liquid water content" ;
		rad_liquid_water:standard_name = "atmosphere_cloud_liquid_water_content" ;
		rad_liquid_water:source = "JMR" ;
		rad_liquid_water:institution = "NASA/JPL" ;
		rad_liquid_water:units = "kg/m^2" ;
		rad_liquid_water:quality_flag = "qual_rad_1hz_tb187 and qual_rad_1hz_tb238 and qual_rad_1hz_tb340 and interp_flag_tb" ;
		rad_liquid_water:scale_factor = 0.01 ;
		rad_liquid_water:coordinates = "lon lat" ;
		rad_liquid_water:comment = "Should not be used over land." ;
	int ice_range_20hz_ku(time, meas_ind) ;
		ice_range_20hz_ku:_FillValue = 2147483647 ;
		ice_range_20hz_ku:long_name = "20 Hz Ku band altimeter range (ice retracking)" ;
		ice_range_20hz_ku:standard_name = "altimeter_range" ;
		ice_range_20hz_ku:units = "m" ;
		ice_range_20hz_ku:add_offset = 1300000. ;
		ice_range_20hz_ku:scale_factor = 0.0001 ;
		ice_range_20hz_ku:coordinates = "lon_20hz lat_20hz" ;
		ice_range_20hz_ku:comment = "Distance antenna-COG (cog_corr), USO drift correction (uso_corr) and internal path correction (internal_path_delay_corr_ku) included" ;
	int ice_range_20hz_c(time, meas_ind) ;
		ice_range_20hz_c:_FillValue = 2147483647 ;
		ice_range_20hz_c:long_name = "20 Hz C band altimeter range (ice retracking)" ;
		ice_range_20hz_c:standard_name = "altimeter_range" ;
		ice_range_20hz_c:units = "m" ;
		ice_range_20hz_c:add_offset = 1300000. ;
		ice_range_20hz_c:scale_factor = 0.0001 ;
		ice_range_20hz_c:coordinates = "lon_20hz lat_20hz" ;
		ice_range_20hz_c:comment = "Distance antenna-COG (cog_corr), USO drift correction (uso_corr) and internal path correction (internal_path_delay_corr_c) included" ;
	short ice_sig0_20hz_ku(time, meas_ind) ;
		ice_sig0_20hz_ku:_FillValue = 32767s ;
		ice_sig0_20hz_ku:long_name = "20 Hz Ku band backscatter coefficient (ice retracking)" ;
		ice_sig0_20hz_ku:standard_name = "surface_backwards_scattering_coefficient_of_radar_wave" ;
		ice_sig0_20hz_ku:units = "dB" ;
		ice_sig0_20hz_ku:scale_factor = 0.01 ;
		ice_sig0_20hz_ku:coordinates = "lon_20hz lat_20hz" ;
		ice_sig0_20hz_ku:comment = "AGC instrumental errors correction and internal calibration correction (internal_corr_sig0_ku) included" ;
	short ice_sig0_20hz_c(time, meas_ind) ;
		ice_sig0_20hz_c:_FillValue = 32767s ;
		ice_sig0_20hz_c:long_name = "20 Hz C band backscatter coefficient (ice retracking)" ;
		ice_sig0_20hz_c:standard_name = "surface_backwards_scattering_coefficient_of_radar_wave" ;
		ice_sig0_20hz_c:units = "dB" ;
		ice_sig0_20hz_c:scale_factor = 0.01 ;
		ice_sig0_20hz_c:coordinates = "lon_20hz lat_20hz" ;
		ice_sig0_20hz_c:comment = "AGC instrumental errors correction and internal calibration correction (internal_corr_sig0_c) included" ;
	byte ice_qual_flag_20hz_ku(time, meas_ind) ;
		ice_qual_flag_20hz_ku:_FillValue = 127b ;
		ice_qual_flag_20hz_ku:long_name = "20 Hz Ku band ice retracking quality flag" ;
		ice_qual_flag_20hz_ku:flag_values = 0b, 1b ;
		ice_qual_flag_20hz_ku:flag_meanings = "good bad" ;
		ice_qual_flag_20hz_ku:coordinates = "lon_20hz lat_20hz" ;
		ice_qual_flag_20hz_ku:comment = "ice retracking quality flag" ;
	short mqe_20hz_ku(time, meas_ind) ;
		mqe_20hz_ku:_FillValue = 32767s ;
		mqe_20hz_ku:long_name = "20 Hz Ku band MQE (ocean retracking)" ;
		mqe_20hz_ku:units = "count" ;
		mqe_20hz_ku:scale_factor = 0.0001 ;
		mqe_20hz_ku:coordinates = "lon_20hz lat_20hz" ;
		mqe_20hz_ku:comment = "Mean Quadratic Error between the waveforms samples and the corresponding model samples built from the ocean retracking outputs" ;
	short mqe_20hz_c(time, meas_ind) ;
		mqe_20hz_c:_FillValue = 32767s ;
		mqe_20hz_c:long_name = "20 Hz C band MQE (ocean retracking)" ;
		mqe_20hz_c:units = "count" ;
		mqe_20hz_c:scale_factor = 0.0001 ;
		mqe_20hz_c:coordinates = "lon_20hz lat_20hz" ;
		mqe_20hz_c:comment = "Mean Quadratic Error between the waveforms samples and the corresponding model samples built from the ocean retracking outputs" ;
	short peakiness_20hz_ku(time, meas_ind) ;
		peakiness_20hz_ku:_FillValue = 32767s ;
		peakiness_20hz_ku:long_name = "20 Hz peakiness on Ku band waveforms" ;
		peakiness_20hz_ku:units = "count" ;
		peakiness_20hz_ku:scale_factor = 0.001 ;
		peakiness_20hz_ku:coordinates = "lon_20hz lat_20hz" ;
	short peakiness_20hz_c(time, meas_ind) ;
		peakiness_20hz_c:_FillValue = 32767s ;
		peakiness_20hz_c:long_name = "20 Hz peakiness on C band waveforms" ;
		peakiness_20hz_c:units = "count" ;
		peakiness_20hz_c:scale_factor = 0.001 ;
		peakiness_20hz_c:coordinates = "lon_20hz lat_20hz" ;
	short ssha(time) ;
		ssha:_FillValue = 32767s ;
		ssha:long_name = "sea surface height anomaly" ;
		ssha:standard_name = "sea_surface_height_above_sea_level" ;
		ssha:source = "Poseidon-2" ;
		ssha:institution = "CNES" ;
		ssha:units = "m" ;
		ssha:scale_factor = 0.001 ;
		ssha:coordinates = "lon lat" ;
		ssha:comment = "= altitude of satellite (alt) - Ku band corrected altimeter range (range_ku) - altimeter ionospheric correction on Ku band (iono_corr_alt_ku) - model dry tropospheric correction (model_dry_tropo_corr) - radiometer wet tropospheric correction (rad_wet_tropo_corr) - sea state bias correction in Ku band (sea_state_bias_ku) - solid earth tide height (solid_earth_tide) - geocentric ocean tide height solution 1 (ocean_tide_sol1) - geocentric pole tide height (pole_tide) - inverted barometer height correction (inv_bar_corr) - high frequency fluctuations of the sea surface topography (hf_fluctuations_corr for I/GDR off line products only) - mean sea surface (mean_sea_surface). Set to default if the altimeter surface type (surface_type) is set to 1, 2, or 3 (lake_enclosed_sea, ice, or land)" ;

// global attributes:
		:Conventions = "CF-1.1" ;
		:title = "GDR - Native dataset" ;
		:institution = "CNES and JPL" ;
		:source = "radar altimeter" ;
		:history = "2016-01-20 14:02:12 : Creation" ;
		:contact = "CNES aviso@altimetry.fr NASA/JPL podaac@podaac.jpl.nasa.gov" ;
		:references = "CNES Reprocessing Tool 2.0 (Updates to time tags, ranges, models and all JMR derived parameters updated with dedicated recalibration of JMR in 2015)" ;
		:processing_center = "SALP and JSDS" ;
		:reference_document = "AVISO and PODAAC User Handbook IGDR and GDR Jason Products, SALP-MU-M5-OP-13184-CN" ;
		:mission_name = "Jason-1" ;
		:altimeter_sensor_name = "POSEIDON-2" ;
		:radiometer_sensor_name = "JMR" ;
		:doris_sensor_name = "2GM" ;
		:gpsr_sensor_name = "TRSR" ;
		:acq_station_name = "CNES/NASA" ;
		:cycle_number = 73 ;
		:absolute_rev_number = 9151 ;
		:pass_number = 13 ;
		:absolute_pass_number = 18301 ;
		:equator_time = "2003-12-30 15:07:28.902000" ;
		:equator_longitude = 289.84 ;
		:first_meas_time = "2003-12-30 14:39:22.759345" ;
		:last_meas_time = "2003-12-30 15:35:34.135558" ;
		:ellipsoid_axis = 6378136.3 ;
		:ellipsoid_flattening = 0.0033528131778969 ;
}
