netcdf CSU_SSMI_FCDR_V01R00_F13_D20030101_S0033_E0215_R40107 {
dimensions:
	npixel_lores = 64 ;
	npixel_hires = 128 ;
	nscan_lores = 1607 ;
	nscan_hires = 3214 ;
	ntest = 9 ;
	numchar = 23 ;
variables:
	double orbit_lores(nscan_lores) ;
		orbit_lores:_FillValue = -9999.9 ;
		orbit_lores:valid_range = 1., 32767. ;
		orbit_lores:long_name = "Fractional orbit number" ;
	double scan_time_lores(nscan_lores) ;
		scan_time_lores:units = "seconds since 1987-01-01T00:00:00.00Z" ;
		scan_time_lores:_FillValue = -9999.9 ;
		scan_time_lores:valid_range = 0., 2000000000. ;
		scan_time_lores:standard_name = "time" ;
		scan_time_lores:long_name = "Scan start time (UTC) for low resolution scans in a referenced or elapsed time format" ;
	char scan_datetime_lores(nscan_lores, numchar) ;
		scan_datetime_lores:_FillValue = "0" ;
		scan_datetime_lores:long_name = "Scan start time (UTC) for low resolution scans in ISO8601 date/time (YYYY-MM-DDTHH-MM-SS.SSZ) format" ;
	float spacecraft_lat_lores(nscan_lores) ;
		spacecraft_lat_lores:units = "degrees_north" ;
		spacecraft_lat_lores:_FillValue = -9999.9f ;
		spacecraft_lat_lores:valid_range = -90.f, 90.f ;
		spacecraft_lat_lores:long_name = "Spacecraft latitude corresponding to scan_time_lores" ;
	float spacecraft_lon_lores(nscan_lores) ;
		spacecraft_lon_lores:units = "degrees_east" ;
		spacecraft_lon_lores:_FillValue = -9999.9f ;
		spacecraft_lon_lores:valid_range = -180.f, 180.f ;
		spacecraft_lon_lores:long_name = "Spacecraft longitude corresponding to scan_time_lores" ;
	float spacecraft_alt_lores(nscan_lores) ;
		spacecraft_alt_lores:units = "km" ;
		spacecraft_alt_lores:_FillValue = -9999.9f ;
		spacecraft_alt_lores:valid_range = 0.f, 1000.f ;
		spacecraft_alt_lores:long_name = "Spacecraft altitude corresponding to scan_time_lores" ;
	float lat_lores(nscan_lores, npixel_lores) ;
		lat_lores:units = "degrees_north" ;
		lat_lores:_FillValue = -9999.9f ;
		lat_lores:valid_range = -90.f, 90.f ;
		lat_lores:standard_name = "latitude" ;
		lat_lores:long_name = "Latitude for low resolution channels" ;
	float lon_lores(nscan_lores, npixel_lores) ;
		lon_lores:units = "degrees_east" ;
		lon_lores:_FillValue = -9999.9f ;
		lon_lores:valid_range = -180.f, 180.f ;
		lon_lores:standard_name = "longitude" ;
		lon_lores:long_name = "Longitude for low resolution channels" ;
	float fcdr_tb19v(nscan_lores, npixel_lores) ;
		fcdr_tb19v:units = "kelvin" ;
		fcdr_tb19v:_FillValue = -9999.9f ;
		fcdr_tb19v:valid_range = 50.f, 350.f ;
		fcdr_tb19v:standard_name = "brightness_temperature" ;
		fcdr_tb19v:long_name = "NOAA FCDR of 19.35 GHz vertically-polarized brightness temperature" ;
		fcdr_tb19v:coordinates = "lon_lores lat_lores" ;
		fcdr_tb19v:grid_mapping = "crs" ;
		fcdr_tb19v:comment = "Calibration Offset applied to 19v channel =  0.00 K (Adjusted to F13)" ;
	float fcdr_tb19h(nscan_lores, npixel_lores) ;
		fcdr_tb19h:units = "kelvin" ;
		fcdr_tb19h:_FillValue = -9999.9f ;
		fcdr_tb19h:valid_range = 50.f, 350.f ;
		fcdr_tb19h:standard_name = "brightness_temperature" ;
		fcdr_tb19h:long_name = "NOAA FCDR of 19.35 GHz horizontally-polarized brightness temperature" ;
		fcdr_tb19h:coordinates = "lon_lores lat_lores" ;
		fcdr_tb19h:grid_mapping = "crs" ;
		fcdr_tb19h:comment = "Calibration Offset applied to 19h channel =  0.00 K (Adjusted to F13)" ;
	float fcdr_tb22v(nscan_lores, npixel_lores) ;
		fcdr_tb22v:units = "kelvin" ;
		fcdr_tb22v:_FillValue = -9999.9f ;
		fcdr_tb22v:valid_range = 50.f, 350.f ;
		fcdr_tb22v:standard_name = "brightness_temperature" ;
		fcdr_tb22v:long_name = "NOAA FCDR of 22.235 GHz vertically-polarized brightness temperature" ;
		fcdr_tb22v:coordinates = "lon_lores lat_lores" ;
		fcdr_tb22v:grid_mapping = "crs" ;
		fcdr_tb22v:comment = "Calibration Offset applied to 22v channel =  0.00 K (Adjusted to F13)" ;
	float fcdr_tb37v(nscan_lores, npixel_lores) ;
		fcdr_tb37v:units = "kelvin" ;
		fcdr_tb37v:_FillValue = -9999.9f ;
		fcdr_tb37v:valid_range = 50.f, 350.f ;
		fcdr_tb37v:standard_name = "brightness_temperature" ;
		fcdr_tb37v:long_name = "NOAA FCDR of 37.0 GHz vertically-polarized brightness temperature" ;
		fcdr_tb37v:coordinates = "lon_lores lat_lores" ;
		fcdr_tb37v:grid_mapping = "crs" ;
		fcdr_tb37v:comment = "Calibration Offset applied to 37v channel =  0.00 K (Adjusted to F13)" ;
	float fcdr_tb37h(nscan_lores, npixel_lores) ;
		fcdr_tb37h:units = "kelvin" ;
		fcdr_tb37h:_FillValue = -9999.9f ;
		fcdr_tb37h:valid_range = 50.f, 350.f ;
		fcdr_tb37h:standard_name = "brightness_temperature" ;
		fcdr_tb37h:long_name = "NOAA FCDR of 37.0 GHz horizontally-polarized brightness temperature" ;
		fcdr_tb37h:coordinates = "lon_lores lat_lores" ;
		fcdr_tb37h:grid_mapping = "crs" ;
		fcdr_tb37h:comment = "Calibration Offset applied to 37h channel =  0.00 K (Adjusted to F13)" ;
	float eia_lores(nscan_lores, npixel_lores) ;
		eia_lores:units = "degrees" ;
		eia_lores:_FillValue = -9999.9f ;
		eia_lores:valid_range = 0.f, 90.f ;
		eia_lores:long_name = "Earth Incidence Angle for low resolution channels" ;
		eia_lores:coordinates = "lon_lores lat_lores" ;
	byte sun_glint_lores(nscan_lores, npixel_lores) ;
		sun_glint_lores:units = "degrees" ;
		sun_glint_lores:_FillValue = -99b ;
		sun_glint_lores:valid_range = -90b, 127b ;
		sun_glint_lores:long_name = "Sun Glint Angle for low resolution channels" ;
		sun_glint_lores:coordinates = "lon_lores lat_lores" ;
	byte quality_lores(nscan_lores, npixel_lores) ;
		quality_lores:valid_range = 0UB, 255UB ;
		quality_lores:long_name = "Quality Flag for low resolution channels" ;
		quality_lores:coordinates = "lon_lores lat_lores" ;
		quality_lores:flag_values = 0b, 1b, 2b, 3b, 4b, 5b, 6b, 7b, 8b, 9b, 10b, 11b, 12b, 13b, 14b, 100b, 101b, 102b, 103b, 104b, 105b, 106b, 107b, 108b, 109b, 110b, 111b, 112b, 113b, 114b, 115b, 116b, 117b, 118b, 119b, 120b, 0b ;
		quality_lores:flag_meanings = "Good_data Possible_sun_glint Climatology_check_warning_(19V_Channel) Climatology_check_warning_(19H_Channel) Climatology_check_warning_(22V_Channel) Climatology_check_warning_(37V_Channel) Climatology_check_warning_(37H_Channel) Climatology_check_warning_(85V_Channel) Climatology_check_warning_(85H_Channel) Climatology_check_warning_(Multiple_low-res_channels) Climatology_check_warning_(Multiple_high-res_channels) Warning adjacent/cross-pol_pixel_flagged_as_bad Warning_of_increased_noise_in_85V_channel_on_DMSP_F08 RADCAL_correction_applied_to_Tb22v_(do_not_use_for_climate) Ta correction made by eliminating spikes in scan cal data Correction made to Ta by correcting for spikes in warm/cold load cal data Data_is_missing_from_file_or_unreadable Geolocation_check_flagged_in_input_BASE_file Climatology_check_flagged_in_input_BASE_file Climatology_check_failed_(19V_Channel) Climatology_check_failed_(19H_Channel) Climatology_check_failed_(22V_Channel) Climatology_check_failed_(37V_Channel) Climatology_check_failed_(37H_Channel) Climatology_check_failed_(85V_Channel) Climatology_check_failed_(85H_Channel) Climatology_check_failed_(Multiple_low-res_channels) Climatology_check_failed_(Multiple_high-res_channels) Distance between pixels is nonphysical Antenna_temperatures_are_<50_or_>350 Lat/Lon_values are_out_of_range Failure_of_85V_channel_on_DMSP_F08 Failure_of_85V_and_increased_noise_in_85H_on_DMSP_F08 Failure_of_both_85V_and_85H_channels_on_DMSP_F08 Invalid_scan_time Ta set to missing due to bad cal data All data set to missing " ;
		quality_lores:comment = "0=Good data, 1-99=Minor issue (use with caution), 100-255=Major issue (set to missing); FLAG VALUES: [0] Good data; [1] Possible sun glint; [2] Climatology check warning (19V Channel); [3] Climatology check warning (19H Channel); [4] Climatology check warning (22V Channel); [5] Climatology check warning (37V Channel); [6] Climatology check warning (37H Channel); [7] Climatology check warning (85V Channel); [8] Climatology check warning (85H Channel); [9] Climatology check warning (Multiple low-res channels); [10] Climatology check warning (Multiple high-res channels); [11] Warning adjacent/cross-pol pixel flagged as bad; [12] Warning of increased noise in 85V channel on DMSP F08; [13] RADCAL correction applied to Tb22v (do not use for climate); [14] Correction made to Ta by correcting for spikes in warm/cold load cal data; [100] Data is missing from file or unreadable; [101] Geolocation check flagged in input BASE file; [102] Climatology check flagged in input BASE file; [103] Climatology check failed (19V Channel); [104] Climatology check failed (19H Channel); [105] Climatology check failed (22V Channel); [106] Climatology check failed (37V Channel); [107] Climatology check failed (37H Channel); [108] Climatology check failed (85V Channel); [109] Climatology check failed (85H Channel); [110] Climatology check failed (Multiple low-res channels); [111] Climatology check failed (Multiple high-res channels); [112] Distance between pixels is nonphysical; [113] Antenna temperatures are < 50 or > 350; [114] Lat/Lon values are out of range; [115] Failure of 85V channel on DMSP F08; [116] Failure of 85V and increased noise in 85H on DMSP F08; [117] Failure of both 85V and 85H channels on DMSP F08; [118] Invalid scan time; [119] Ta set to missing due to bad cal data; [120] All data set to missing; " ;
	double orbit_hires(nscan_hires) ;
		orbit_hires:_FillValue = -9999.9 ;
		orbit_hires:valid_range = 1., 32767. ;
		orbit_hires:long_name = "Fractional orbit number" ;
	double scan_time_hires(nscan_hires) ;
		scan_time_hires:units = "seconds since 1987-01-01T00:00:00.00Z" ;
		scan_time_hires:_FillValue = -9999.9 ;
		scan_time_hires:valid_range = 0., 2000000000. ;
		scan_time_hires:standard_name = "time" ;
		scan_time_hires:long_name = "Scan start time (UTC) for high resolution scans in a referenced or elapsed time format" ;
	char scan_datetime_hires(nscan_hires, numchar) ;
		scan_datetime_hires:_FillValue = "0" ;
		scan_datetime_hires:long_name = "Scan start time (UTC) for high resolution scans in ISO8601 date/time (YYYY-MM-DDTHH-MM-SS.SSZ) format" ;
	float spacecraft_lat_hires(nscan_hires) ;
		spacecraft_lat_hires:units = "degrees_north" ;
		spacecraft_lat_hires:_FillValue = -9999.9f ;
		spacecraft_lat_hires:valid_range = -90.f, 90.f ;
		spacecraft_lat_hires:long_name = "Spacecraft latitude corresponding to scan_time_hires" ;
	float spacecraft_lon_hires(nscan_hires) ;
		spacecraft_lon_hires:units = "degrees_east" ;
		spacecraft_lon_hires:_FillValue = -9999.9f ;
		spacecraft_lon_hires:valid_range = -180.f, 180.f ;
		spacecraft_lon_hires:long_name = "Spacecraft longitude corresponding to scan_time_hires" ;
	float spacecraft_alt_hires(nscan_hires) ;
		spacecraft_alt_hires:units = "km" ;
		spacecraft_alt_hires:_FillValue = -9999.9f ;
		spacecraft_alt_hires:valid_range = 0.f, 1000.f ;
		spacecraft_alt_hires:long_name = "Spacecraft altitude corresponding to scan_time_hires" ;
	float lat_hires(nscan_hires, npixel_hires) ;
		lat_hires:units = "degrees_north" ;
		lat_hires:_FillValue = -9999.9f ;
		lat_hires:valid_range = -90.f, 90.f ;
		lat_hires:standard_name = "latitude" ;
		lat_hires:long_name = "Latitude for high resolution channels" ;
	float lon_hires(nscan_hires, npixel_hires) ;
		lon_hires:units = "degrees_east" ;
		lon_hires:_FillValue = -9999.9f ;
		lon_hires:valid_range = -180.f, 180.f ;
		lon_hires:standard_name = "longitude" ;
		lon_hires:long_name = "Longitude for high resolution channels" ;
	float fcdr_tb85v(nscan_hires, npixel_hires) ;
		fcdr_tb85v:units = "kelvin" ;
		fcdr_tb85v:_FillValue = -9999.9f ;
		fcdr_tb85v:valid_range = 50.f, 350.f ;
		fcdr_tb85v:standard_name = "brightness_temperature" ;
		fcdr_tb85v:long_name = "NOAA FCDR of 85.5 GHz vertically-polarized brightness temperature" ;
		fcdr_tb85v:coordinates = "lon_hires lat_hires" ;
		fcdr_tb85v:grid_mapping = "crs" ;
		fcdr_tb85v:comment = "Calibration Offset applied to 85v channel =  0.00 K (Adjusted to F13)" ;
	float fcdr_tb85h(nscan_hires, npixel_hires) ;
		fcdr_tb85h:units = "kelvin" ;
		fcdr_tb85h:_FillValue = -9999.9f ;
		fcdr_tb85h:valid_range = 50.f, 350.f ;
		fcdr_tb85h:standard_name = "brightness_temperature" ;
		fcdr_tb85h:long_name = "NOAA FCDR of 85.5 GHz horizontally-polarized brightness temperature" ;
		fcdr_tb85h:coordinates = "lon_hires lat_hires" ;
		fcdr_tb85h:grid_mapping = "crs" ;
		fcdr_tb85h:comment = "Calibration Offset applied to 85h channel =  0.00 K (Adjusted to F13)" ;
	float eia_hires(nscan_hires, npixel_hires) ;
		eia_hires:units = "degrees" ;
		eia_hires:_FillValue = -9999.9f ;
		eia_hires:valid_range = 0.f, 90.f ;
		eia_hires:long_name = "Earth Incidence Angle for high resolution channels" ;
		eia_hires:coordinates = "lon_hires lat_hires" ;
	byte sun_glint_hires(nscan_hires, npixel_hires) ;
		sun_glint_hires:units = "degrees" ;
		sun_glint_hires:_FillValue = -99b ;
		sun_glint_hires:valid_range = -90b, 127b ;
		sun_glint_hires:long_name = "Sun Glint Angle for high resolution channels" ;
		sun_glint_hires:coordinates = "lon_hires lat_hires" ;
	byte quality_hires(nscan_hires, npixel_hires) ;
		quality_hires:valid_range = 0UB, 255UB ;
		quality_hires:long_name = "Quality Flag for high resolution channels" ;
		quality_hires:coordinates = "lon_hires lat_hires" ;
		quality_hires:flag_values = 0b, 1b, 2b, 3b, 4b, 5b, 6b, 7b, 8b, 9b, 10b, 11b, 12b, 13b, 14b, 100b, 101b, 102b, 103b, 104b, 105b, 106b, 107b, 108b, 109b, 110b, 111b, 112b, 113b, 114b, 115b, 116b, 117b, 118b, 119b, 120b, 0b ;
		quality_hires:flag_meanings = "Good_data Possible_sun_glint Climatology_check_warning_(19V_Channel) Climatology_check_warning_(19H_Channel) Climatology_check_warning_(22V_Channel) Climatology_check_warning_(37V_Channel) Climatology_check_warning_(37H_Channel) Climatology_check_warning_(85V_Channel) Climatology_check_warning_(85H_Channel) Climatology_check_warning_(Multiple_low-res_channels) Climatology_check_warning_(Multiple_high-res_channels) Warning adjacent/cross-pol_pixel_flagged_as_bad Warning_of_increased_noise_in_85V_channel_on_DMSP_F08 RADCAL_correction_applied_to_Tb22v_(do_not_use_for_climate) Ta correction made by eliminating spikes in scan cal data Correction made to Ta by correcting for spikes in warm/cold load cal data Data_is_missing_from_file_or_unreadable Geolocation_check_flagged_in_input_BASE_file Climatology_check_flagged_in_input_BASE_file Climatology_check_failed_(19V_Channel) Climatology_check_failed_(19H_Channel) Climatology_check_failed_(22V_Channel) Climatology_check_failed_(37V_Channel) Climatology_check_failed_(37H_Channel) Climatology_check_failed_(85V_Channel) Climatology_check_failed_(85H_Channel) Climatology_check_failed_(Multiple_low-res_channels) Climatology_check_failed_(Multiple_high-res_channels) Distance between pixels is nonphysical Antenna_temperatures_are_<50_or_>350 Lat/Lon_values are_out_of_range Failure_of_85V_channel_on_DMSP_F08 Failure_of_85V_and_increased_noise_in_85H_on_DMSP_F08 Failure_of_both_85V_and_85H_channels_on_DMSP_F08 Invalid_scan_time Ta set to missing due to bad cal data All data set to missing " ;
		quality_hires:comment = "0=Good data, 1-99=Minor issue (use with caution), 100-255=Major issue (set to missing); FLAG VALUES: [0] Good data; [1] Possible sun glint; [2] Climatology check warning (19V Channel); [3] Climatology check warning (19H Channel); [4] Climatology check warning (22V Channel); [5] Climatology check warning (37V Channel); [6] Climatology check warning (37H Channel); [7] Climatology check warning (85V Channel); [8] Climatology check warning (85H Channel); [9] Climatology check warning (Multiple low-res channels); [10] Climatology check warning (Multiple high-res channels); [11] Warning adjacent/cross-pol pixel flagged as bad; [12] Warning of increased noise in 85V channel on DMSP F08; [13] RADCAL correction applied to Tb22v (do not use for climate); [14] Correction made to Ta by correcting for spikes in warm/cold load cal data; [100] Data is missing from file or unreadable; [101] Geolocation check flagged in input BASE file; [102] Climatology check flagged in input BASE file; [103] Climatology check failed (19V Channel); [104] Climatology check failed (19H Channel); [105] Climatology check failed (22V Channel); [106] Climatology check failed (37V Channel); [107] Climatology check failed (37H Channel); [108] Climatology check failed (85V Channel); [109] Climatology check failed (85H Channel); [110] Climatology check failed (Multiple low-res channels); [111] Climatology check failed (Multiple high-res channels); [112] Distance between pixels is nonphysical; [113] Antenna temperatures are < 50 or > 350; [114] Lat/Lon values are out of range; [115] Failure of 85V channel on DMSP F08; [116] Failure of 85V and increased noise in 85H on DMSP F08; [117] Failure of both 85V and 85H channels on DMSP F08; [118] Invalid scan time; [119] Ta set to missing due to bad cal data; [120] All data set to missing; " ;
	int quality_tests(ntest) ;
		quality_tests:long_name = "Results from quality control tests" ;
		quality_tests:flag_values = 1b, 2b, 3b, 4b, 5b, 6b, 7b, 8b, 9b ;
		quality_tests:flag_meanings = "Number_of_nonphysical_or_bad_pixel_values Number_of_pixels_with_bad_geolocation Number_of_scans_with_geolocation_error_in_input_BASE_file Number_of_scans_with_climatology_error_in_input_BASE_file Number_of_scans_corrected_for_calibration/temperature_spike Number_of_scans_flagged_missing_due_to_calibration/temperature_spike Number_of_scans_with_errors_in_geolocation Number_of_scans_with_sensor_errors Number_of_scans_exceeding_specified_variance_from_climatological_values " ;
		quality_tests:comment = "Results from quality control tests; Test 1: Number of nonphysical or bad pixel values; Test 2: Number of pixels with bad geolocation; Test 3: Number of scans with geolocation error in input BASE file; Test 4: Number of scans with climatology error in input BASE file; Test 5: Number of scans corrected for calibration/temperature spike; Test 6: Number of scans flagged missing due to calibration/temperature spike; Test 7: Number of scans with errors in geolocation; Test 8: Number of scans with sensor errors; Test 9: Number of scans exceeding specified variance from climatological values; " ;
	float nominal_elevation_angle ;
		nominal_elevation_angle:units = "degrees" ;
		nominal_elevation_angle:valid_range = 0.f, 90.f ;
		nominal_elevation_angle:long_name = "Nominal sensor elevation angle" ;
	float delta_elevation_angle ;
		delta_elevation_angle:units = "degrees" ;
		delta_elevation_angle:valid_range = -2.f, 2.f ;
		delta_elevation_angle:long_name = "Offset in the sensor elevation angle from nominal" ;
	float spacecraft_roll ;
		spacecraft_roll:units = "degrees" ;
		spacecraft_roll:valid_range = -2.f, 2.f ;
		spacecraft_roll:standard_name = "platform_roll_angle" ;
		spacecraft_roll:long_name = "Spacecraft roll angle offset from nominal" ;
	float spacecraft_pitch ;
		spacecraft_pitch:units = "degrees" ;
		spacecraft_pitch:valid_range = -2.f, 2.f ;
		spacecraft_pitch:standard_name = "platform_pitch_angle" ;
		spacecraft_pitch:long_name = "Spacecraft pitch angle offset from nominal" ;
	float spacecraft_yaw ;
		spacecraft_yaw:units = "degrees" ;
		spacecraft_yaw:valid_range = -2.f, 2.f ;
		spacecraft_yaw:standard_name = "platform_yaw_angle" ;
		spacecraft_yaw:long_name = "Spacecraft yaw angle offset from nominal" ;
	char crs ;
		crs:long_name = "coordinate reference system" ;
		crs:grid_mapping_name = "latitude_longitude" ;
		crs:longitude_of_prime_meridian = 0.f ;
		crs:semi_major_axis = 6378.14f ;
		crs:semi_minor_axis = 6356.755f ;
		crs:mean_earth_radius = 6371.f ;
		crs:inverse_flattening = 298.2572f ;

// global attributes:
		:Conventions = "CF-1.6" ;
		:Metadata_Conventions = "CF-1.6, Unidata Dataset Discovery v1.0, NOAA CDR v1.0, GDS v2.0" ;
		:standard_name_vocabulary = "CF Standard Name Table (v20, 11 September 2012)" ;
		:id = "CSU_SSMI_FCDR_V01R00_F13_D20030101_S0033_E0215_R40107.nc" ;
		:naming_authority = "gov.noaa.ncdc" ;
		:metadata_link = "gov.noaa.ncdc:C00827" ;
		:title = "CSU SSM/I FCDR" ;
		:product_version = "V01R00" ;
		:revision_date = "2013-02-01" ;
		:summary = "Colorado State University Special Sensor Microwave/Imager (SSM/I) Fundamental Climate Data Record (FCDR) of intercalibrated brightness temperatures" ;
		:keywords = "EARTH SCIENCE > SPECTRAL/ENGINEERING > MICROWAVE > BRIGHTNESS TEMPERATURE" ;
		:keywords_vocabulary = "NASA Global Change Master Directory (GCMD) Earth Science Keywords, Version 6.0" ;
		:platform = "DMSP 5D-2/F13 > Defense Meteorological Satellite Program-F13" ;
		:sensor = "SSM/I > Special Sensor Microwave/Imager" ;
		:cdm_data_type = "Swath" ;
		:cdr_program = "NOAA Climate Data Record Program for satellites, FY 2013" ;
		:cdr_variable = "fcdr_tb19v, fcdr_tb19h, fcdr_tb22v, fcdr_tb37v, fcdr_tb37h, fcdr_tb85v, fcdr_tb85h" ;
		:source = "SSMI_TDRBASE_V01R03_F13_D20030101_S0033_E0215_R40107.nc" ;
		:date_created = "2013-02-02T22:28MST" ;
		:creator_name = "Wesley Berg" ;
		:creator_url = "http://rain.atmos.colostate.edu/FCDR" ;
		:creator_email = "fcdr@atmos.colostate.edu" ;
		:institution = "Colorado State University, Dept. of Atmospheric Science, Kummerow research group" ;
		:processing_level = "NOAA Level 2" ;
		:geospatial_lat_min = " -87.78" ;
		:geospatial_lat_max = "  87.52" ;
		:geospatial_lon_min = "-180.00" ;
		:geospatial_lon_max = " 180.00" ;
		:geospatial_lat_units = "degrees_north" ;
		:geospatial_lon_units = "degrees_east" ;
		:spatial_resolution = "19 V/H GHz: 43km X 69km, 22 V GHz: 40km X 50km, 37 V/H GHz: 28km X 37km, 85 V/H GHz: 13km X 15km" ;
		:time_coverage_start = "2003-01-01T00:33:32Z" ;
		:time_coverage_end = "2003-01-01T02:15:23Z" ;
		:time_coverage_duration = "PT1H41M51S" ;
		:license = "No restrictions on access or use" ;
		:contributor_name = "Christian Kummerow, Wesley Berg, Mathew Sapiano" ;
		:contributor_role = "Principal investigator, Co-Investigator and developer with overall responsibility for FCDR data software and documentation, Responsible for intercalibration geolocation and cross-track bias adjustments including associated software and documentation" ;
		:orbit_number = "40107" ;
}
