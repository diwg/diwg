netcdf S5P_TEST_L1B_RA_BD6_20140827T114200_20140827T115800_53811_01_000901_20141209T120000 {

// global attributes:
		:Conventions = "CF-1.6" ;
		:institution = "KNMI" ;
		:library_information = "\n../lib/libCOREFoundation.so (TROPOMI L01b CORE library) v0.9.1.14380 Build 201511162052 by tropdev@bhltrdev.knmi.nl\n../lib/libGeo.so (TROPOMI L01b Geolocation library) v0.9.1.14380 Build 201511162053 by tropdev@bhltrdev.knmi.nl\n../lib/libMath.so (TROPOMI L01b MATH library) v0.9.1.14380 Build 201511162053 by tropdev@bhltrdev.knmi.nl\n../lib/TROP_L0InputSubsystem.so (TROPOMI L0 Input Subsystem) v0.9.1 Build Nov 17 2015 07:49:59\n../lib/TROP_KeyDataSubSystem.so (TROPOMI Key Data Input Subsystem) v0.9.1 Build Nov 17 2015 07:50:28\n../lib/TROP_L1BOutputSubsystem.so (TROPOMI L1b Output Subsystem) v0.9.1 Build Nov 17 2015 07:50:27" ;
		:orbit = 53811 ;
		:processor_version = "0.9.1.14380_local" ;
		:summary = "Radiance product band 6 (NIR detector)" ;
		:time_coverage_end = "2014-08-27T11:51:47Z" ;
		:time_coverage_start = "2014-08-27T11:45:53Z" ;
		:time_reference = "2014-08-27T00:00:00Z" ;
		:title = "Sentinel-5p TROPOMI Level 1b Radiance product band 6 (NIR detector)" ;

group: BAND6_RADIANCE {

  group: STANDARD_MODE {
    dimensions:
    	time = 1 ;
    	scanline = 326 ; // flight direction
    	spectral_channel = 497 ; // spectral dimension
    	ground_pixel = 448 ; // scan direction (perpendicular to flight direction)
    	ncorner = 4 ;
    	nsettings = 5 ;
    	nbinningregions = 18 ;

    group: OBSERVATIONS {
      types:
        float(*) vlen_float ;
      variables:
      	int scanline(scanline) ;
      		scanline:comment = "This dimension variable defines the indices along track; index starts at 0" ;
      		scanline:long_name = "along track dimension index" ;
      		scanline:units = "1" ;
      	int delta_time(time, scanline) ;
      		delta_time:comment = "Time difference with time for each measurement" ;
      		delta_time:_FillValue = -2147483647 ;
      		delta_time:long_name = "offset from the reference start time of measurement" ;
      		delta_time:units = "milliseconds since 2014-08-27 00:00:00" ;
      	int spectral_channel(spectral_channel) ;
      		spectral_channel:comment = "This dimension variable defines the indices spectral dimension; index starts at 0" ;
      		spectral_channel:long_name = "wavelength dimension index" ;
      		spectral_channel:units = "1" ;
      	ushort detector_column_qualification(time, scanline, spectral_channel) ;
      		detector_column_qualification:comment = "Qualification flag indicating column indicating column type or state" ;
      		detector_column_qualification:units = "1" ;
      		detector_column_qualification:_FillValue = 65535US ;
      		detector_column_qualification:flag_values = 0US, 1US, 16US, 32US, 64US, 256US, 512US, 1024US, 2048US ;
      		detector_column_qualification:flag_masks = 0US, 1US, 16US, 98US, 98US, 3840US, 3840US, 3840US, 3840US ;
      		detector_column_qualification:flag_meanings = "no_qualification skipped uvn_odd uvn_prepost uvn_overscan swir_adc0 swir_adc1 swir_adc2 swir_adc3" ;
      		detector_column_qualification:long_name = "Detector column qualification flags" ;
      		detector_column_qualification:max_val = 65534US ;
      		detector_column_qualification:min_val = 0US ;
      	int ground_pixel(ground_pixel) ;
      		ground_pixel:comment = "This dimension variable defines the indices across track; index starts at 0" ;
      		ground_pixel:long_name = "across track dimension index" ;
      		ground_pixel:units = "1" ;
      	ushort detector_row_qualification(time, scanline, ground_pixel) ;
      		detector_row_qualification:comment = "Qualification flag indicating row type or state" ;
      		detector_row_qualification:_FillValue = 65535US ;
      		detector_row_qualification:flag_values = 0US, 1US, 2US, 4US, 8US, 16US, 256US, 4096US, 8192US ;
      		detector_row_qualification:flag_masks = 0US, 9US, 2US, 4US, 9US, 16US, 256US, 4096US, 8192US ;
      		detector_row_qualification:flag_meanings = "no_qualification uvn_ror uvn_dump uvn_covered uvn_overscan uvn_higain swir_reference gen_transistion gen_non_illuminated" ;
      		detector_row_qualification:long_name = "Detector row qualification flags" ;
      		detector_row_qualification:max_val = 65534US ;
      		detector_row_qualification:min_val = 0US ;
      		detector_row_qualification:units = "1" ;
      	ubyte ground_pixel_quality(time, scanline, ground_pixel) ;
      		ground_pixel_quality:comment = "Quality assessment information for each ground pixel" ;
      		ground_pixel_quality:coordinates = "longitude latitude" ;
      		ground_pixel_quality:max_val = 254UB ;
      		ground_pixel_quality:_FillValue = 255UB ;
      		ground_pixel_quality:flag_values = 0UB, 1UB, 2UB, 4UB, 8UB, 16UB, 128UB ;
      		ground_pixel_quality:flag_masks = 0UB, 1UB, 2UB, 4UB, 8UB, 16UB, 128UB ;
      		ground_pixel_quality:flag_meanings = "no_error solar_eclipse sun_glint_possible descending night geo_boundary_crossing geolocation_error" ;
      		ground_pixel_quality:long_name = "ground pixel quality flag" ;
      		ground_pixel_quality:min_val = 0UB ;
      		ground_pixel_quality:units = "1" ;
      	ushort measurement_quality(time, scanline) ;
      		measurement_quality:flag_masks = 0US, 1US, 2US, 16US, 32US, 128US, 256US, 4096US ;
      		measurement_quality:flag_meanings = "no_error proc_skipped no_residual saa spacecraft_manoeuvre sub_grp irr_out_of_range sub_group" ;
      		measurement_quality:long_name = "measurement quality flag" ;
      		measurement_quality:max_val = 65534US ;
      		measurement_quality:min_val = 0US ;
      		measurement_quality:units = "1" ;
      		measurement_quality:comment = "Overall quality information for a measurement" ;
      		measurement_quality:coordinates = "longitude latitude" ;
      		measurement_quality:_FillValue = 65535US ;
      		measurement_quality:flag_values = 0US, 1US, 2US, 16US, 32US, 128US, 256US, 4096US ;
      	ubyte quality_level(time, scanline, ground_pixel, spectral_channel) ;
      		quality_level:comment = "Overall quality assessment information for each (spectral) pixel" ;
      		quality_level:coordinates = "longitude latitude" ;
      		quality_level:_FillValue = 255UB ;
      		quality_level:long_name = "qualiy level of spectral channel" ;
      		quality_level:max_val = 100UB ;
      		quality_level:min_val = 0UB ;
      		quality_level:units = "1" ;
      	float radiance(time, scanline, ground_pixel, spectral_channel) ;
      		radiance:ancilary_vars = "radiance_noise radiance_error quality_level spectral_channel_quality ground_pixel_quality" ;
      		radiance:coordinates = "longitude latitude" ;
      		radiance:comment = "Measured spectral radiance for each spectral pixel" ;
      		radiance:_FillValue = 9.96921e+36f ;
      		radiance:long_name = "spectral photon radiance" ;
      		radiance:units = "mol.m-2.nm-1.sr-1.s-1" ;
      	byte radiance_error(time, scanline, ground_pixel, spectral_channel) ;
      		radiance_error:comment = "The radiance_error is a measure for the one standard deviation error of the bias of the radiance measurement; it is expressed in decibel (dB), i.e. 10 times the base-10 logarithmic value of the ratio between the radiance and the estimation error." ;
      		radiance_error:coordinates = "longitude latitude" ;
      		radiance_error:_FillValue = -127b ;
      		radiance_error:long_name = "spectral photon radiance error, one standard deviation" ;
      		radiance_error:units = "1" ;
      	byte radiance_noise(time, scanline, ground_pixel, spectral_channel) ;
      		radiance_noise:coordinates = "longitude latitude" ;
      		radiance_noise:comment = "The radiance_noise is a measure for the one standard deviation random error of the radiance measurement; it is expressed in decibel (dB), i.e. 10 times the base-10 logarithmic value of the ratio between the radiance and the random error." ;
      		radiance_noise:_FillValue = -127b ;
      		radiance_noise:long_name = "spectral photon radiance noise, one standard deviation" ;
      		radiance_noise:units = "1" ;
      	vlen_float small_pixel_radiance(time, scanline, ground_pixel) ;
      		small_pixel_radiance:long_name = "small pixel photon radiance" ;
      		small_pixel_radiance:units = "mol.m-2.nm-1.sr-1.s-1" ;
      		small_pixel_radiance:comment = "Measured spectral radiance for the spectral channel dedicated for the small pixel measurements" ;
      		small_pixel_radiance:coordinates = "longitude latitude" ;
      	ubyte spectral_channel_quality(time, scanline, ground_pixel, spectral_channel) ;
      		spectral_channel_quality:comment = "Quality assessment information for each (spectral) pixel" ;
      		spectral_channel_quality:units = "1" ;
      		spectral_channel_quality:coordinates = "longitude latitude" ;
      		spectral_channel_quality:_FillValue = 255UB ;
      		spectral_channel_quality:flag_values = 0UB, 1UB, 2UB, 8UB, 16UB, 32UB, 64UB, 128UB ;
      		spectral_channel_quality:flag_masks = 0UB, 1UB, 2UB, 8UB, 16UB, 32UB, 64UB, 128UB ;
      		spectral_channel_quality:flag_meanings = "no_error missing bad_pixel processing_error saturated transient rts underflow" ;
      		spectral_channel_quality:long_name = "spectral channel quality flag" ;
      		spectral_channel_quality:max_val = 254UB ;
      		spectral_channel_quality:min_val = 0UB ;
      	int time(time) ;
      		time:comment = "Reference time of the measurements. The reference time is set to yyyy-mm-ddT00:00:00 UTC, where yyyy-mm-dd is the day on which the measurements of a particular data granule start." ;
      		time:long_name = "reference start time of measurement" ;
      		time:standard_name = "time" ;
      		time:units = "seconds since 2010-01-01 00:00:00" ;
      } // group OBSERVATIONS

    group: GEODATA {
      variables:
      	float earth_sun_distance(time) ;
      		earth_sun_distance:comment = "1 ua equals 149,597,870,700 meters" ;
      		earth_sun_distance:_FillValue = 9.96921e+36f ;
      		earth_sun_distance:units = "ua" ;
      		earth_sun_distance:long_name = "distance between the earth and the sun" ;
      		earth_sun_distance:max_val = 1.02f ;
      		earth_sun_distance:min_val = 0.98f ;
      	float latitude_bounds(time, scanline, ground_pixel, ncorner) ;
      		latitude_bounds:comment = "The four latitude boundaries of each ground pixel." ;
      		latitude_bounds:_FillValue = 9.96921e+36f ;
      		latitude_bounds:units = "degrees north" ;
      	float latitude(time, scanline, ground_pixel) ;
      		latitude:comment = "Latitude of the center of each ground pixel on the WGS84  reference ellipsoid" ;
      		latitude:_FillValue = 9.96921e+36f ;
      		latitude:long_name = "pixel center latitude" ;
      		latitude:max_val = 90.f ;
      		latitude:min_val = -90.f ;
      		latitude:standard_name = "latitude" ;
      		latitude:bounds = "latitude_bounds" ;
      		latitude:units = "degrees north" ;
      	float longitude_bounds(time, scanline, ground_pixel, ncorner) ;
      		longitude_bounds:comment = "The four longitude boundaries of each ground pixel." ;
      		longitude_bounds:_FillValue = 9.96921e+36f ;
      		longitude_bounds:units = "degrees east" ;
      	float longitude(time, scanline, ground_pixel) ;
      		longitude:comment = "Longitude of the center of each ground pixel on the WGS84 reference ellipsoid" ;
      		longitude:_FillValue = 9.96921e+36f ;
      		longitude:long_name = "pixel center longitude" ;
      		longitude:bounds = "longitude_bounds" ;
      		longitude:max_val = 180.f ;
      		longitude:min_val = -180.f ;
      		longitude:standard_name = "longitude" ;
      		longitude:units = "degrees east" ;
      	float satellite_altitude(time, scanline) ;
      		satellite_altitude:comment = "The altitude of the spacecraft relative to the WGS84 reference ellipsoid" ;
      		satellite_altitude:_FillValue = 9.96921e+36f ;
      		satellite_altitude:long_name = "satellite altitude" ;
      		satellite_altitude:max_val = 900000.f ;
      		satellite_altitude:min_val = 700000.f ;
      		satellite_altitude:units = "m" ;
      	float satellite_latitude(time, scanline) ;
      		satellite_latitude:comment = "Latitude of the spacecraft sub-satellite point on the WGS84 reference ellipsoid" ;
      		satellite_latitude:_FillValue = 9.96921e+36f ;
      		satellite_latitude:long_name = "sub-satellite latitude" ;
      		satellite_latitude:max_val = 90.f ;
      		satellite_latitude:min_val = -90.f ;
      		satellite_latitude:units = "degrees north" ;
      	float satellite_longitude(time, scanline) ;
      		satellite_longitude:comment = "Longitude of the spacecraft sub-satellite point on the WGS84 reference ellipsoid" ;
      		satellite_longitude:_FillValue = 9.96921e+36f ;
      		satellite_longitude:max_val = 180.f ;
      		satellite_longitude:min_val = -180.f ;
      		satellite_longitude:units = "degrees east" ;
      	float satellite_orbit_phase(time, scanline) ;
      		satellite_orbit_phase:comment = "Relative offset (0.0 ... 1.0) of the measurement in the orbit" ;
      		satellite_orbit_phase:_FillValue = 9.96921e+36f ;
      		satellite_orbit_phase:long_name = "fractional satellite orbit phase" ;
      		satellite_orbit_phase:max_val = 1.02f ;
      		satellite_orbit_phase:min_val = -0.02f ;
      		satellite_orbit_phase:units = "1" ;
      	float solar_azimuth_angle(time, scanline, ground_pixel) ;
      		solar_azimuth_angle:units = "degree" ;
      		solar_azimuth_angle:comment = "Solar azimuth angle at the ground pixel location on the reference ellipsoid. Angle is measured clockwise from the North (East = 90, South = 180, West = 270)" ;
      		solar_azimuth_angle:coordinates = "longitude latitude" ;
      		solar_azimuth_angle:_FillValue = 9.96921e+36f ;
      		solar_azimuth_angle:long_name = "solar azimuth angle" ;
      		solar_azimuth_angle:max_val = 360.f ;
      		solar_azimuth_angle:min_val = 0.f ;
      		solar_azimuth_angle:standard_name = "solar_azimuth_angle" ;
      	float solar_zenith_angle(time, scanline, ground_pixel) ;
      		solar_zenith_angle:comment = "Solar zenith angle at the ground pixel location on the reference ellipsoid. Angle is measured away from the vertical. ESA definition of day side: SZA less the 92 degrees" ;
      		solar_zenith_angle:coordinates = "longitude latitude" ;
      		solar_zenith_angle:_FillValue = 9.96921e+36f ;
      		solar_zenith_angle:long_name = "solar zenith angle" ;
      		solar_zenith_angle:max_val = 180.f ;
      		solar_zenith_angle:min_val = 0.f ;
      		solar_zenith_angle:standard_name = "solar_zenith_angle" ;
      		solar_zenith_angle:units = "degree" ;
      	float viewing_azimuth_angle(time, scanline, ground_pixel) ;
      		viewing_azimuth_angle:comment = "Azimuth angle of the satellite at the ground pixel location on the reference ellipsoid. Angle is measured clockwise from the North (East = 90, South = 180, West = 270)" ;
      		viewing_azimuth_angle:coordinates = "longitude latitude" ;
      		viewing_azimuth_angle:_FillValue = 9.96921e+36f ;
      		viewing_azimuth_angle:units = "degree" ;
      		viewing_azimuth_angle:long_name = "viewing azimuth angle" ;
      		viewing_azimuth_angle:max_val = 360.f ;
      		viewing_azimuth_angle:min_val = 0.f ;
      		viewing_azimuth_angle:standard_name = "platform_azimuth_angle" ;
      	float viewing_zenith_angle(time, scanline, ground_pixel) ;
      		viewing_zenith_angle:comment = "Zenith angle of the satellite at the ground pixel location on the reference ellipsoid. Angle is measured away from the vertical." ;
      		viewing_zenith_angle:coordinates = "longitude latitude" ;
      		viewing_zenith_angle:_FillValue = 9.96921e+36f ;
      		viewing_zenith_angle:long_name = "viewing zenith angle" ;
      		viewing_zenith_angle:max_val = 180.f ;
      		viewing_zenith_angle:min_val = 0.f ;
      		viewing_zenith_angle:standard_name = "platform_zenith_angle" ;
      		viewing_zenith_angle:units = "degree" ;
      } // group GEODATA

    group: INSTRUMENT {
      types:
        compound housekeeping_data_type {
          float temp_det1 ;
          float temp_det2 ;
          float temp_det3 ;
          float temp_det4 ;
          float data_offset_s ;
          float temp_tss_up_neg_x ;
          float temp_tss_up_neg_y ;
          float temp_tss_up_pos_x ;
          float temp_tss_up_pos_y ;
          float temp_tss_up_mid ;
          float temp_tss_low_mid ;
          float temp_low_uvn_obm ;
          float temp_up_uvn_obm ;
          float temp_obm_swir ;
          float temp_obm_solar_baffle ;
          float temp_cu_sls_stim ;
          float temp_obm_swir_grating ;
          float temp_obm_swir_if ;
          float temp_pelt_cu_sls1 ;
          float temp_pelt_cu_sls2 ;
          float temp_pelt_cu_sls3 ;
          float temp_pelt_cu_sls4 ;
          float temp_pelt_cu_sls5 ;
          ubyte difm_status ;
          ubyte fmm_status ;
          ubyte det1_led_status ;
          ubyte det2_led_status ;
          ubyte det3_led_status ;
          ubyte det4_led_status ;
          ubyte common_led_status ;
          ubyte sls1_status ;
          ubyte sls2_status ;
          ubyte sls3_status ;
          ubyte sls4_status ;
          ubyte sls5_status ;
          ubyte wls_status ;
          ubyte filler_char1 ;
          float swir_vdet_bias ;
        }; // housekeeping_data_type
        compound housekeeping_data_type_str {
          string temp_det1 ;
          string temp_det2 ;
          string temp_det3 ;
          string temp_det4 ;
          string data_offset_s ;
          string temp_tss_up_neg_x ;
          string temp_tss_up_neg_y ;
          string temp_tss_up_pos_x ;
          string temp_tss_up_pos_y ;
          string temp_tss_up_mid ;
          string temp_tss_low_mid ;
          string temp_low_uvn_obm ;
          string temp_up_uvn_obm ;
          string temp_obm_swir ;
          string temp_obm_solar_baffle ;
          string temp_cu_sls_stim ;
          string temp_obm_swir_grating ;
          string temp_obm_swir_if ;
          string temp_pelt_cu_sls1 ;
          string temp_pelt_cu_sls2 ;
          string temp_pelt_cu_sls3 ;
          string temp_pelt_cu_sls4 ;
          string temp_pelt_cu_sls5 ;
          string difm_status ;
          string fmm_status ;
          string det1_led_status ;
          string det2_led_status ;
          string det3_led_status ;
          string det4_led_status ;
          string common_led_status ;
          string sls1_status ;
          string sls2_status ;
          string sls3_status ;
          string sls4_status ;
          string sls5_status ;
          string wls_status ;
          string filler_char1 ;
          string swir_vdet_bias ;
        }; // housekeeping_data_type_str
        compound instrument_configuration_type {
          int ic_id ;
          short ic_version ;
        }; // instrument_configuration_type
        compound instrument_configuration_type_str {
          string ic_id ;
          string ic_version ;
        }; // instrument_configuration_type_str
        compound msmt_to_det_row_table_type {
          short det_start_row ;
          short det_end_row ;
        }; // msmt_to_det_row_table_type
        compound msmt_to_det_row_table_type_str {
          string det_start_row ;
          string det_end_row ;
        }; // msmt_to_det_row_table_type_str
        compound binning_table_type {
          short size ;
          short binning_factor ;
          short gain ;
          short detector_start_row ;
          short detector_stop_row ;
          short measurement_start_row ;
          short measurement_stop_row ;
        }; // binning_table_type
        compound binning_table_type_str {
          string size ;
          string binning_factor ;
          string gain ;
          string detector_stop_row ;
          string detector_start_row ;
          string measurement_start_row ;
          string measurement_stop_row ;
        }; // binning_table_type_str
        compound instrument_settings_type {
          int ic_id ;
          short ic_version ;
          short ic_set ;
          short ic_idx ;
          short processing_class ;
          float master_cycle_period ;
          float coaddition_period ;
          float exposure_time ;
          float msmt_mcp_ft_offset ;
          float msmt_ft_msmt_start_offset ;
          float msmt_duration ;
          float flush_duration ;
          short nr_coadditions ;
          short cds_gain ;
          float pga_gain ;
          float dac_offset ;
          int master_cycle_period_us ;
          int coaddition_period_us ;
          int exposure_time_us ;
          int exposure_period_us ;
          short small_pixel_column ;
          short stop_column_read ;
          short start_column_coad ;
          short stop_column_coad ;
          short pga_gain_code ;
          short dac_offset_code ;
          ubyte clock_mode ;
          ubyte clipping ;
        }; // instrument_settings_type
        compound instrument_settings_type_str {
          string ic_id ;
          string ic_version ;
          string ic_set ;
          string ic_idx ;
          string processing_class ;
          string master_cycle_period ;
          string coaddition_period ;
          string exposure_time ;
          string msmt_mcp_ft_offset ;
          string msmt_ft_msmt_start_offset ;
          string msmt_duration ;
          string flush_duration ;
          string nr_coadditions ;
          string cds_gain ;
          string pga_gain ;
          string dac_offset ;
          string master_cycle_period_us ;
          string coaddition_period_us ;
          string exposure_time_us ;
          string exposure_period_us ;
          string pga_gain_code ;
          string dac_offset_code ;
          string small_pixel_column ;
          string stop_column_read ;
          string start_column_coad ;
          string stop_column_coad ;
          string clock_mode ;
          string clipping ;
        }; // instrument_settings_type_str
      variables:
      	housekeeping_data_type housekeeping_data(time, scanline) ;
      		housekeeping_data_type housekeeping_data:_FillValue = 
          {9.96921e+36, 9.96921e+36, 9.96921e+36, 9.96921e+36, 9.96921e+36, 9.96921e+36, 9.96921e+36, 9.96921e+36, 9.96921e+36, 9.96921e+36, 9.96921e+36, 9.96921e+36, 9.96921e+36, 9.96921e+36, 9.96921e+36, 9.96921e+36, 9.96921e+36, 9.96921e+36, 9.96921e+36, 9.96921e+36, 9.96921e+36, 9.96921e+36, 9.96921e+36, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 9.96921e+36} ;
      		housekeeping_data_type_str housekeeping_data:units = 
          {"K", "K", "K", "K", "s", "K", "K", "K", "K", "K", "K", "K", "K", "K", "K", "K", "K", "K", "K", "K", "K", "K", "K", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "V"} ;
      		housekeeping_data:comment = "Fields that describe scanline dependent instrument characteristics, like detector temperatures, etc." ;
      	instrument_configuration_type instrument_configuration(time, scanline) ;
      		instrument_configuration_type instrument_configuration:_FillValue = 
          {-2147483647, -32767} ;
      		instrument_configuration_type_str instrument_configuration:units = {"1", "1"} ;
      		instrument_configuration:long_name = "instrument configuration, IcID and IcVersion" ;
      		instrument_configuration:comment = "The Instrument Configuration ID defines the type of measurement and its purposes. The number of Instrument Configuration IDs will increase over the mission as new types of measurements are created / used; The Instrument Configuration Version allows to differentiate between multiple versions for a specific IcID." ;
      	msmt_to_det_row_table_type measurement_to_detector_row_table(time, scanline, ground_pixel) ;
      		msmt_to_det_row_table_type_str measurement_to_detector_row_table:units = {"1", "1"} ;
      		msmt_to_det_row_table_type measurement_to_detector_row_table:_FillValue = {-32767, -32767} ;
      		measurement_to_detector_row_table:comment = "Conversion table from measurement row to begin and end row on detector" ;
      	float nominal_wavelength(time, ground_pixel, spectral_channel) ;
      		nominal_wavelength:comment = "The nominal spectral wavelength for each cross track pixel as a function of the spectral channel." ;
      		nominal_wavelength:units = "1e-09 m" ;
      		nominal_wavelength:_FillValue = 9.96921e+36f ;
      		nominal_wavelength:long_name = "spectral channel nominal wavelength" ;
      		nominal_wavelength:standard_name = "radiation_wavelength" ;
      	short processing_class(time, scanline) ;
      		processing_class:comment = "The processing_class defines the type of measurement at a very high level. Contrary to Instrument Configuration IDs, only a limited, fixed set of processing classes is identified. Examples of processing classes are Earth_radiance, Sun_irradiance, CLED, WLS, Dark, Background, ...;" ;
      		processing_class:_FillValue = -32767s ;
      		processing_class:long_name = "processing class" ;
      		processing_class:max_val = 255s ;
      		processing_class:min_val = 0s ;
      		processing_class:units = "1" ;
      	int sample_cycle(time, scanline) ;
      		sample_cycle:comment = "sample_cycle provides a sample_cycle index for each scanline; index starts at 0" ;
      		sample_cycle:_FillValue = -2147483647 ;
      		sample_cycle:long_name = "sample cycle" ;
      		sample_cycle:units = "1" ;
      	int sample_cycle_length(time, scanline) ;
      		sample_cycle_length:comment = "Length of sample_cycle" ;
      		sample_cycle_length:_FillValue = -2147483647 ;
      		sample_cycle_length:long_name = "length of sample cycle" ;
      		sample_cycle_length:units = "ms" ;
      	binning_table_type binning_table(nsettings, nbinningregions) ;
      		binning_table_type binning_table:_FillValue = 
          {-32767, -32767, -32767, -32767, -32767, -32767, -32767} ;
      		binning_table_type_str binning_table:units = 
          {"1", "1", "1", "1", "1", "1", "1"} ;
      		binning_table_type_str binning_table:comment = 
          {"Number of rows in the area before binning / read-out", "Binning factor for the area; 0 if rows are skipped", "CCD output gain for the area (0 = dump, 1 = 1x, 2 = 2x)", "Start row of the binning area on the detector", "Stop row of the binning area on the detector; the stop row is exclusive (i.e. up to, but not including)", "Start row of the binning area in the measurement. Set to -1 in case the area is skipped. Reflects the rows that are actually written to the output, in case a subset of the data is written.", "Stop row of the binning area in the measurement; the stop row is exclusive (i.e. up to, but not including). Set to -1 in case the area is skipped. Reflects the rows that are actually written to the output, in case a subset of the data is written."} ;
      		binning_table:long_name = "binning table settings" ;
      	instrument_settings_type instrument_settings(nsettings) ;
      		instrument_settings_type instrument_settings:_FillValue = 
          {-2147483647, -32767, -32767, -32767, -32767, 9.96921e+36, 9.96921e+36, 9.96921e+36, 9.96921e+36, 9.96921e+36, 9.96921e+36, 9.96921e+36, -32767, -32767, 9.96921e+36, 9.96921e+36, -2147483647, -2147483647, -2147483647, -2147483647, -32767, -32767, -32767, -32767, -32767, -32767, 255, 255} ;
      		instrument_settings_type_str instrument_settings:units = 
          {"1", "1", "1", "1", "1", "s", "s", "s", "s", "s", "s", "s", "1", "1", "1", "V", "us", "us", "us", "us", "1", "1", "1", "1", "1", "1", "1", "1"} ;
      		instrument_settings:comment = "All fields that determine the instrument configuration and are relevant for data processing, like exposure tme, binning factors, co-addition period, gain settings, status of calibration unit, etc." ;
      } // group INSTRUMENT
    } // group STANDARD_MODE
  } // group BAND6_RADIANCE

group: METADATA {

  group: ESA_METADATA {

    // group attributes:
    		:objectType = "Earth_Explorer_File" ;

    group: earth_explorer_header {

      // group attributes:
      		:objectType = "Earth_Explorer_Header" ;

      group: fixed_header {

        // group attributes:
        		:File_Class = "OFFL" ;
        		:File_Description = "Sentinel-5p TROPOMI Level 1b Radiance product band 6 (NIR detector)" ;
        		:File_Name = "S5P_TEST_L1B_RA_BD6_20140827T114200_20140827T115800_53811_01_000901_20141209T120000" ;
        		:File_Type = "L1B_RA_BD6" ;
        		:File_Version = "L1B_RA_BD6" ;
        		:Mission = "Sentinel-5P" ;
        		:Notes = " " ;
        		:objectType = "Fixed_Header" ;

        group: source {

          // group attributes:
          		:Creation_Date = "UTC=2015-11-18T08:25:24" ;
          		:Creator = "KNMI TROPOMI L01b processor" ;
          		:Creator_Version = "0.9.1.14380_local" ;
          		:System = "DLR PDGS" ;
          		:objectType = "Source" ;
          } // group source

        group: validity_period {

          // group attributes:
          		:Validity_Start = "UTC=2014-08-27T11:42:00" ;
          		:Validity_Stop = "UTC=2014-08-27T11:58:00" ;
          		:objectType = "Validity_Period" ;
          } // group validity_period
        } // group fixed_header

      group: variable_header {

        // group attributes:
        		:objectType = "Variable_Header" ;

        group: gmd\:lineage {

          // group attributes:
          		:objectType = "gmd:LI_Lineage" ;
          		:gmd\:statement = "L1b  dataset produced by the DLR PDGS from the S5p TROPOMI L0 product" ;

          group: gmd\:processStep {

            // group attributes:
            		:gmd\:description = "Processing of L0 to L1b data using the KNMI TROPOMI L01b processor" ;
            		:objectType = "gmi:LE_ProcessStep" ;

            group: gmd\:source\#09 {

              // group attributes:
              		:gmd\:description = "L0 Band 5 NIR science data" ;
              		:objectType = "gmi:LE_Source" ;

              group: gmi\:processedLevel {

                // group attributes:
                		:gmd\:code = "L0" ;
                		:objectType = "gmd:MD_Identifier" ;
                } // group gmi\:processedLevel

              group: gmd\:sourceCitation {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2015-11-18" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeListValue = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date

                group: gmd\:title {

                  // group attributes:
                  		:gco\:characterString = "L0 instrument data for band 5" ;
                  } // group gmd\:title

                group: gmd\:alternateTitle\#1 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_TEST_L0__ODB_4__20140827T114000_20140827T114500_53811_00.RAW" ;
                  } // group gmd\:alternateTitle\#1

                group: gmd\:alternateTitle\#2 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_TEST_L0__ODB_4__20140827T114500_20140827T115000_53811_01.RAW" ;
                  } // group gmd\:alternateTitle\#2

                group: gmd\:alternateTitle\#3 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_TEST_L0__ODB_4__20140827T115000_20140827T115500_53811_02.RAW" ;
                  } // group gmd\:alternateTitle\#3

                group: gmd\:alternateTitle\#4 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_TEST_L0__ODB_4__20140827T115500_20140827T120000_53811_03.RAW" ;
                  } // group gmd\:alternateTitle\#4
                } // group gmd\:sourceCitation
              } // group gmd\:source\#09

            group: gmd\:source\#08 {

              // group attributes:
              		:gmd\:description = "L0 Band 4 VIS science data" ;
              		:objectType = "gmi:LE_Source" ;

              group: gmi\:processedLevel {

                // group attributes:
                		:gmd\:code = "L0" ;
                		:objectType = "gmd:MD_Identifier" ;
                } // group gmi\:processedLevel

              group: gmd\:sourceCitation {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2015-11-18" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeListValue = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date

                group: gmd\:title {

                  // group attributes:
                  		:gco\:characterString = "L0 instrument data for band 4" ;
                  } // group gmd\:title

                group: gmd\:alternateTitle\#1 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_TEST_L0__ODB_3__20140827T114000_20140827T114500_53811_00.RAW" ;
                  } // group gmd\:alternateTitle\#1

                group: gmd\:alternateTitle\#2 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_TEST_L0__ODB_3__20140827T114500_20140827T115000_53811_01.RAW" ;
                  } // group gmd\:alternateTitle\#2

                group: gmd\:alternateTitle\#3 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_TEST_L0__ODB_3__20140827T115000_20140827T115500_53811_02.RAW" ;
                  } // group gmd\:alternateTitle\#3

                group: gmd\:alternateTitle\#4 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_TEST_L0__ODB_3__20140827T115500_20140827T120000_53811_03.RAW" ;
                  } // group gmd\:alternateTitle\#4
                } // group gmd\:sourceCitation
              } // group gmd\:source\#08

            group: gmd\:source\#11 {

              // group attributes:
              		:gmd\:description = "L0 Band 7 SWIR science data" ;
              		:objectType = "gmi:LE_Source" ;

              group: gmi\:processedLevel {

                // group attributes:
                		:gmd\:code = "L0" ;
                		:objectType = "gmd:MD_Identifier" ;
                } // group gmi\:processedLevel

              group: gmd\:sourceCitation {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2015-11-18" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeListValue = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date

                group: gmd\:title {

                  // group attributes:
                  		:gco\:characterString = "L0 instrument data for band 7" ;
                  } // group gmd\:title

                group: gmd\:alternateTitle\#1 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_TEST_L0__ODB_6__20140827T114000_20140827T114500_53811_00.RAW" ;
                  } // group gmd\:alternateTitle\#1

                group: gmd\:alternateTitle\#2 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_TEST_L0__ODB_6__20140827T114500_20140827T115000_53811_01.RAW" ;
                  } // group gmd\:alternateTitle\#2

                group: gmd\:alternateTitle\#3 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_TEST_L0__ODB_6__20140827T115000_20140827T115500_53811_02.RAW" ;
                  } // group gmd\:alternateTitle\#3

                group: gmd\:alternateTitle\#4 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_TEST_L0__ODB_6__20140827T115500_20140827T120000_53811_03.RAW" ;
                  } // group gmd\:alternateTitle\#4
                } // group gmd\:sourceCitation
              } // group gmd\:source\#11

            group: gmd\:source\#01 {

              // group attributes:
              		:gmd\:description = "Auxiliary Calibration Key Data product" ;
              		:objectType = "gmi:LE_Source" ;

              group: gmd\:sourceCitation {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2015-11-18" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeListValue = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date

                group: gmd\:title {

                  // group attributes:
                  		:gco\:characterString = "Auxiliary Calibration Key Data Set" ;
                  } // group gmd\:title

                group: gmd\:alternateTitle\#1 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_TEST_AUX_L1_CKD_20140101T000000_20151231T000000_00000_01_000900_20150915T120000.h5" ;
                  } // group gmd\:alternateTitle\#1
                } // group gmd\:sourceCitation
              } // group gmd\:source\#01

            group: gmd\:source\#13 {

              // group attributes:
              		:gmd\:description = "L0 Ancillary data" ;
              		:objectType = "gmi:LE_Source" ;

              group: gmi\:processedLevel {

                // group attributes:
                		:gmd\:code = "L0" ;
                		:objectType = "gmd:MD_Identifier" ;
                } // group gmi\:processedLevel

              group: gmd\:sourceCitation {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2015-11-18" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeListValue = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date

                group: gmd\:title {

                  // group attributes:
                  		:gco\:characterString = "L0 instrument ancillary data" ;
                  } // group gmd\:title

                group: gmd\:alternateTitle\#1 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_TEST_L0__SAT_A__20140827T114000_20140827T114500_53811_00.RAW" ;
                  } // group gmd\:alternateTitle\#1

                group: gmd\:alternateTitle\#2 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_TEST_L0__SAT_A__20140827T114500_20140827T115000_53811_01.RAW" ;
                  } // group gmd\:alternateTitle\#2

                group: gmd\:alternateTitle\#3 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_TEST_L0__SAT_A__20140827T115000_20140827T115500_53811_02.RAW" ;
                  } // group gmd\:alternateTitle\#3

                group: gmd\:alternateTitle\#4 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_TEST_L0__SAT_A__20140827T115500_20140827T120000_53811_03.RAW" ;
                  } // group gmd\:alternateTitle\#4
                } // group gmd\:sourceCitation
              } // group gmd\:source\#13

            group: gmd\:source\#03 {

              group: gmd\:sourceCitation {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2015-11-18" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeListValue = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date

                group: gmd\:title {

                  // group attributes:
                  		:gco\:characterString = "In-flight Calibration Key Data Set UVN" ;
                  } // group gmd\:title

                group: gmd\:alternateTitle\#1 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_TEST_ICM_CKDSIR_20140101T000000_20151231T000000_00000_01_000900_20150915T120000.h5" ;
                  } // group gmd\:alternateTitle\#1
                } // group gmd\:sourceCitation
              } // group gmd\:source\#03

            group: gmd\:source\#02 {

              // group attributes:
              		:gmd\:description = "In-flight UVN Calibration Key Data product" ;
              		:objectType = "gmi:LE_Source" ;

              group: gmd\:sourceCitation {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2015-11-18" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeListValue = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date

                group: gmd\:title {

                  // group attributes:
                  		:gco\:characterString = "In-flight Calibration Key Data Set UVN" ;
                  } // group gmd\:title

                group: gmd\:alternateTitle\#1 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_TEST_ICM_CKDUVN_20140101T000000_20151231T000000_00000_01_000900_20150915T120000.h5" ;
                  } // group gmd\:alternateTitle\#1
                } // group gmd\:sourceCitation
              } // group gmd\:source\#02

            group: gmd\:source\#05 {

              // group attributes:
              		:gmd\:description = "L0 Band 1 UV science data" ;
              		:objectType = "gmi:LE_Source" ;

              group: gmi\:processedLevel {

                // group attributes:
                		:gmd\:code = "L0" ;
                		:objectType = "gmd:MD_Identifier" ;
                } // group gmi\:processedLevel

              group: gmd\:sourceCitation {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2015-11-18" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeListValue = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date

                group: gmd\:title {

                  // group attributes:
                  		:gco\:characterString = "L0 instrument data for band 1" ;
                  } // group gmd\:title

                group: gmd\:alternateTitle\#1 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_TEST_L0__ODB_8__20140827T114000_20140827T114500_53811_00.RAW" ;
                  } // group gmd\:alternateTitle\#1

                group: gmd\:alternateTitle\#2 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_TEST_L0__ODB_8__20140827T114500_20140827T115000_53811_01.RAW" ;
                  } // group gmd\:alternateTitle\#2

                group: gmd\:alternateTitle\#3 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_TEST_L0__ODB_8__20140827T115000_20140827T115500_53811_02.RAW" ;
                  } // group gmd\:alternateTitle\#3

                group: gmd\:alternateTitle\#4 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_TEST_L0__ODB_8__20140827T115500_20140827T120000_53811_03.RAW" ;
                  } // group gmd\:alternateTitle\#4
                } // group gmd\:sourceCitation
              } // group gmd\:source\#05

            group: gmd\:source\#04 {

              // group attributes:
              		:gmd\:description = "L0 Engineering data" ;
              		:objectType = "gmi:LE_Source" ;

              group: gmi\:processedLevel {

                // group attributes:
                		:gmd\:code = "L0" ;
                		:objectType = "gmd:MD_Identifier" ;
                } // group gmi\:processedLevel

              group: gmd\:sourceCitation {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2015-11-18" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeListValue = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date

                group: gmd\:title {

                  // group attributes:
                  		:gco\:characterString = "L0 instrument engineering data" ;
                  } // group gmd\:title

                group: gmd\:alternateTitle\#1 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_TEST_L0__ENG_A__20140827T114000_20140827T114500_53811_00.RAW" ;
                  } // group gmd\:alternateTitle\#1

                group: gmd\:alternateTitle\#2 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_TEST_L0__ENG_A__20140827T114500_20140827T115000_53811_01.RAW" ;
                  } // group gmd\:alternateTitle\#2

                group: gmd\:alternateTitle\#3 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_TEST_L0__ENG_A__20140827T115000_20140827T115500_53811_02.RAW" ;
                  } // group gmd\:alternateTitle\#3

                group: gmd\:alternateTitle\#4 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_TEST_L0__ENG_A__20140827T115500_20140827T120000_53811_03.RAW" ;
                  } // group gmd\:alternateTitle\#4
                } // group gmd\:sourceCitation
              } // group gmd\:source\#04

            group: gmd\:source\#07 {

              // group attributes:
              		:gmd\:description = "L0 Band 3 VIS science data" ;
              		:objectType = "gmi:LE_Source" ;

              group: gmi\:processedLevel {

                // group attributes:
                		:gmd\:code = "L0" ;
                		:objectType = "gmd:MD_Identifier" ;
                } // group gmi\:processedLevel

              group: gmd\:sourceCitation {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2015-11-18" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeListValue = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date

                group: gmd\:title {

                  // group attributes:
                  		:gco\:characterString = "L0 instrument data for band 3" ;
                  } // group gmd\:title

                group: gmd\:alternateTitle\#1 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_TEST_L0__ODB_2__20140827T114000_20140827T114500_53811_00.RAW" ;
                  } // group gmd\:alternateTitle\#1

                group: gmd\:alternateTitle\#2 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_TEST_L0__ODB_2__20140827T114500_20140827T115000_53811_01.RAW" ;
                  } // group gmd\:alternateTitle\#2

                group: gmd\:alternateTitle\#3 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_TEST_L0__ODB_2__20140827T115000_20140827T115500_53811_02.RAW" ;
                  } // group gmd\:alternateTitle\#3

                group: gmd\:alternateTitle\#4 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_TEST_L0__ODB_2__20140827T115500_20140827T120000_53811_03.RAW" ;
                  } // group gmd\:alternateTitle\#4
                } // group gmd\:sourceCitation
              } // group gmd\:source\#07

            group: gmd\:source\#06 {

              // group attributes:
              		:gmd\:description = "L0 Band 2 UV science data" ;
              		:objectType = "gmi:LE_Source" ;

              group: gmi\:processedLevel {

                // group attributes:
                		:gmd\:code = "L0" ;
                		:objectType = "gmd:MD_Identifier" ;
                } // group gmi\:processedLevel

              group: gmd\:sourceCitation {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2015-11-18" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeListValue = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date

                group: gmd\:title {

                  // group attributes:
                  		:gco\:characterString = "L0 instrument data for band 2" ;
                  } // group gmd\:title

                group: gmd\:alternateTitle\#1 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_TEST_L0__ODB_1__20140827T114000_20140827T114500_53811_00.RAW" ;
                  } // group gmd\:alternateTitle\#1

                group: gmd\:alternateTitle\#2 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_TEST_L0__ODB_1__20140827T114500_20140827T115000_53811_01.RAW" ;
                  } // group gmd\:alternateTitle\#2

                group: gmd\:alternateTitle\#3 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_TEST_L0__ODB_1__20140827T115000_20140827T115500_53811_02.RAW" ;
                  } // group gmd\:alternateTitle\#3

                group: gmd\:alternateTitle\#4 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_TEST_L0__ODB_1__20140827T115500_20140827T120000_53811_03.RAW" ;
                  } // group gmd\:alternateTitle\#4
                } // group gmd\:sourceCitation
              } // group gmd\:source\#06

            group: gmd\:source\#12 {

              // group attributes:
              		:gmd\:description = "L0 Band 8 SWIR science data" ;
              		:objectType = "gmi:LE_Source" ;

              group: gmi\:processedLevel {

                // group attributes:
                		:gmd\:code = "L0" ;
                		:objectType = "gmd:MD_Identifier" ;
                } // group gmi\:processedLevel

              group: gmd\:sourceCitation {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2015-11-18" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeListValue = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date

                group: gmd\:title {

                  // group attributes:
                  		:gco\:characterString = "L0 instrument data for band 8" ;
                  } // group gmd\:title

                group: gmd\:alternateTitle\#1 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_TEST_L0__ODB_7__20140827T114000_20140827T114500_53811_00.RAW" ;
                  } // group gmd\:alternateTitle\#1

                group: gmd\:alternateTitle\#2 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_TEST_L0__ODB_7__20140827T114500_20140827T115000_53811_01.RAW" ;
                  } // group gmd\:alternateTitle\#2

                group: gmd\:alternateTitle\#3 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_TEST_L0__ODB_7__20140827T115000_20140827T115500_53811_02.RAW" ;
                  } // group gmd\:alternateTitle\#3

                group: gmd\:alternateTitle\#4 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_TEST_L0__ODB_7__20140827T115500_20140827T120000_53811_03.RAW" ;
                  } // group gmd\:alternateTitle\#4
                } // group gmd\:sourceCitation
              } // group gmd\:source\#12

            group: gmi\:report {

              // group attributes:
              		:gmi\:description = "L0 processed to L1b data using the KNMI TROPOMI L01b processor" ;
              		:gmi\:fileType = "netCDF" ;
              		:gmi\:name = "TROPOMI L01b processing report" ;
              		:objectType = "gmi:LE_ProcessStepReport" ;
              } // group gmi\:report

            group: gmi\:processingInformation {

              // group attributes:
              		:objectType = "gmi:LE_Processing" ;

              group: gmi\:softwareReference {

                // group attributes:
                		:gmd\:title = "L01b processor description" ;
                		:objectType = "gmd:CI_Citation" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2014-12-31" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeListValue = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date
                } // group gmi\:softwareReference

              group: gmi\:documentation\#1 {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;
                		:gmd\:title = "S5P-KNMI-L01B-0009-SD-algorithm_theoretical_basis_document-3.0.0-20140707.pdf" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2014-07-07" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeListValue = "publication" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date
                } // group gmi\:documentation\#1

              group: gmi\:identifier {

                // group attributes:
                		:gmd\:code = "KNMI TROPOMI L01b processor" ;
                		:objectType = "gmd:MD_Identifier" ;
                } // group gmi\:identifier

              group: gmi\:documentation\#2 {

                // group attributes:
                		:gmd\:title = "S5P-KNMI-L01B-0012-SD-input_output_data_specification-3.0.0-20140707.pdf" ;
                		:objectType = "gmd:CI_Citation" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2014-07-07" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeListValue = "publication" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date
                } // group gmi\:documentation\#2
              } // group gmi\:processingInformation

            group: gmi\:output {

              // group attributes:
              		:gmd\:description = "TROPOMI L1b Radiance product band 6 (NIR detector)" ;
              		:objectType = "gmi:LE_Source" ;

              group: gmi\:processedLevel {

                // group attributes:
                		:gmd\:code = "L1b" ;
                		:objectType = "gmd:MD_Identifier" ;
                } // group gmi\:processedLevel

              group: gmd\:sourceCitation {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;
                		:gmd\:title = "S5P_TEST_L1B_RA_BD6_20140827T114200_20140827T115800_53811_01_000901_20141209T120000" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2015-11-18" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeListValue = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date
                } // group gmd\:sourceCitation
              } // group gmi\:output

            group: gmd\:source\#10 {

              // group attributes:
              		:gmd\:description = "L0 Band 6 NIR science data" ;
              		:objectType = "gmi:LE_Source" ;

              group: gmi\:processedLevel {

                // group attributes:
                		:gmd\:code = "L0" ;
                		:objectType = "gmd:MD_Identifier" ;
                } // group gmi\:processedLevel

              group: gmd\:sourceCitation {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2015-11-18" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeListValue = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date

                group: gmd\:title {

                  // group attributes:
                  		:gco\:characterString = "L0 instrument data for band 6" ;
                  } // group gmd\:title

                group: gmd\:alternateTitle\#1 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_TEST_L0__ODB_5__20140827T114000_20140827T114500_53811_00.RAW" ;
                  } // group gmd\:alternateTitle\#1

                group: gmd\:alternateTitle\#2 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_TEST_L0__ODB_5__20140827T114500_20140827T115000_53811_01.RAW" ;
                  } // group gmd\:alternateTitle\#2

                group: gmd\:alternateTitle\#3 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_TEST_L0__ODB_5__20140827T115000_20140827T115500_53811_02.RAW" ;
                  } // group gmd\:alternateTitle\#3

                group: gmd\:alternateTitle\#4 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_TEST_L0__ODB_5__20140827T115500_20140827T120000_53811_03.RAW" ;
                  } // group gmd\:alternateTitle\#4
                } // group gmd\:sourceCitation
              } // group gmd\:source\#10
            } // group gmd\:processStep
          } // group gmd\:lineage
        } // group variable_header
      } // group earth_explorer_header
    } // group ESA_METADATA

  group: EOP_METADATA {

    // group attributes:
    		:gml\:id = "S5P_TEST_L1B_RA_BD6_20140827T114200_20140827T115800_53811_01_000901_20141209T120000.EO" ;
    		:objectType = "atm:EarthObservation" ;

    group: eop\:metaDataProperty {

      // group attributes:
      		:eop\:acquisitionType = "NOMINAL" ;
      		:eop\:identifier = "S5P_TEST_L1B_RA_BD6_20140827T114200_20140827T115800_53811_01_000901_20141209T120000" ;
      		:eop\:parentIdentifier = "urn:ogc:def:EOP:ESA:SENTINEL.S5P_TROP_L1B_RA_BD6" ;
      		:eop\:productType = "S5P_OPER_L1B_RA_BD6" ;
      		:eop\:status = "ACQUIRED" ;
      		:objectType = "eop:EarthObservationMetaData" ;

      group: eop\:processing {

        // group attributes:
        		:eop\:nativeProductFormat = "netCDF" ;
        		:eop\:processingCenter = "DLR-DFD" ;
        		:eop\:processingDate = "20151118082524Z" ;
        		:eop\:processingLevel = "L1b" ;
        		:eop\:processorName = "tropl01b" ;
        		:eop\:processorVersion = "0.9.1.14380_local" ;
        		:objectType = "eop:ProcessingInformation" ;
        } // group eop\:processing
      } // group eop\:metaDataProperty

    group: om\:phenomenonTime {

      // group attributes:
      		:gml\:beginPosition = "2014-08-27T11:45:53Z" ;
      		:gml\:endPosition = "2014-08-27T11:51:47Z" ;
      		:objectType = "gml:TimePeriod" ;
      } // group om\:phenomenonTime

    group: om\:featureOfInterest {

      // group attributes:
      		:objectType = "eop:Footprint" ;
      		:gml\:id = "S5P_TEST_L1B_RA_BD6_20140827T114200_20140827T115800_53811_01_000901_20141209T120000.FP" ;

      group: eop\:multiExtentOf {

        // group attributes:
        		:objectType = "gml:MultiSurface" ;

        group: gml\:surfaceMembers {

          // group attributes:
          		:objectType = "gml:Polygon" ;
          		:srsName = "urn:ogc:def:crs:EPSG::4326" ;

          group: gml\:exterior {

            // group attributes:
            		:gml\:posList = "NULL" ;
            		:objectType = "gml:LinearRing" ;
            } // group gml\:exterior
          } // group gml\:surfaceMembers
        } // group eop\:multiExtentOf
      } // group om\:featureOfInterest

    group: om\:observedProperty {

      // group attributes:
      		:nilReason = "inapplicable" ;
      } // group om\:observedProperty

    group: om\:procedure {

      // group attributes:
      		:gml\:id = "S5P_TEST_L1B_RA_BD6_20140827T114200_20140827T115800_53811_01_000901_20141209T120000.EOE" ;
      		:objectType = "eop:EarthObservationEquipment" ;

      group: eop\:instrument {

        // group attributes:
        		:eop\:shortName = "TROPOMI" ;
        		:objectType = "eop:Instrument" ;
        } // group eop\:instrument

      group: eop\:platform {

        // group attributes:
        		:eop\:shortName = "Sentinel-5p" ;
        		:objectType = "eop:Platform" ;
        } // group eop\:platform

      group: eop\:sensor {

        // group attributes:
        		:eop\:sensorType = "ATMOSPHERIC" ;
        		:objectType = "eop:Sensor" ;
        } // group eop\:sensor

      group: eop\:acquisitionParameters {

        // group attributes:
        		:eop\:orbitNumber = "53811" ;
        		:objectType = "eop:Acquisition" ;
        } // group eop\:acquisitionParameters
      } // group om\:procedure
    } // group EOP_METADATA

  group: ISO_METADATA {

    // group attributes:
    		:gmd\:dateStamp = "2015-11-18" ;
    		:gmd\:fileIdentifier = "../data/output/S5P_TEST_L1B_RA_BD6_20140827T114200_20140827T115800_53811_01_000901_20141209T12000.xml" ;
    		:gmd\:metadataStandardName = "ISO 19115-2 Geographic Information - Metadata Part 2 Extensions for imagery and gridded data" ;
    		:gmd\:metadataStandardVersion = "ISO 19115-2:2009(E), S5P profile" ;
    		:objectType = "gmi:MI_Metadata" ;

    group: gmi\:acquisitionInformation {

      // group attributes:
      		:objectType = "gmi:MI_AcquisitionInformation" ;

      group: gmi\:platform {

        // group attributes:
        		:gmi\:description = "Sentinel 5 Precursor" ;
        		:objectType = "gmi:MI_Platform" ;

        group: gmi\:instrument {

          // group attributes:
          		:objectType = "gmi:MI_Instrument" ;

          group: gmi\:type {

            // group attributes:
            		:codeList = " " ;
            		:codeListValue = "UV-VIS-NIR-SWIR imaging spectrometer" ;
            		:objectType = "gmd:MI_SensorTypeCode" ;
            } // group gmi\:type

          group: gmi\:identifier {

            // group attributes:
            		:gmd\:code = "TROPOMI" ;
            		:gmd\:codeSpace = "http://www.esa.int/" ;
            		:objectType = "gmd:RS_Identifier" ;
            } // group gmi\:identifier
          } // group gmi\:instrument

        group: gmi\:identifier {

          // group attributes:
          		:gmd\:code = "S5p" ;
          		:gmd\:codeSpace = "http://www.esa.int/" ;
          		:objectType = "gmd:RS_Identifier" ;
          } // group gmi\:identifier
        } // group gmi\:platform
      } // group gmi\:acquisitionInformation

    group: gmd\:hierarchyLevel {

      // group attributes:
      		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#MD_ScopeCode" ;
      		:codeListValue = "dataset" ;
      		:objectType = "gmd:MD_ScopeCode" ;
      } // group gmd\:hierarchyLevel

    group: gmd\:identificationInfo {

      // group attributes:
      		:gmd\:abstract = "S5p TROPOMI instrument measures..." ;
      		:gmd\:credit = "Financial support by NSO" ;
      		:gmd\:language = "eng" ;
      		:gmd\:topicCategory = "climatologyMeteorologyAtmosphere" ;
      		:objectType = "gmd:MD_DataIdentification" ;

      group: gmd\:citation {

        // group attributes:
        		:gmd\:title = "S5p TROPOMI L1b Radiance product band 6 (NIR detector)" ;
        		:objectType = "gmd:CI_Citation" ;

        group: gmd\:date {

          // group attributes:
          		:gmd\:date = "2015-11-18" ;
          		:objectType = "gmd:CI_Date" ;

          group: gmd\:dateType {

            // group attributes:
            		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
            		:codeListValue = "creation" ;
            		:objectType = "gmd:CI_DateTypeCode" ;
            } // group gmd\:dateType
          } // group gmd\:date

        group: gmd\:identifier {

          // group attributes:
          		:gmd\:code = "../data/output/S5P_TEST_L1B_RA_BD6_20140827T114200_20140827T115800_53811_01_000901_20141209T12000" ;
          		:objectType = "gmd:MD_Identifier" ;
          } // group gmd\:identifier
        } // group gmd\:citation

      group: gmd\:resourceConstraints {

        // group attributes:
        		:gmd\:useLimitation = "no conditions apply" ;
        		:objectType = "gmd:MD_LegalConstraints" ;

        group: gmd\:accessConstraints {

          // group attributes:
          		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#MD_RestrictionCode" ;
          		:codeListValue = "copyright" ;
          		:objectType = "gmd:MD_RestrictionCode" ;
          } // group gmd\:accessConstraints
        } // group gmd\:resourceConstraints

      group: gmd\:extent {

        // group attributes:
        		:objectType = "gmd:EX_Extent" ;

        group: gmd\:temporalElement {

          // group attributes:
          		:objectType = "gmd:EX_TemporalExtent" ;

          group: gmd\:extent {

            // group attributes:
            		:gml\:beginPosition = "2014-08-27T11:45:53Z" ;
            		:gml\:endPosition = "2014-08-27T11:51:47Z" ;
            		:objectType = "gml:TimePeriod" ;
            } // group gmd\:extent
          } // group gmd\:temporalElement

        group: gmd\:geographicElement {

          // group attributes:
          		:extentTypeCode = "true" ;
          		:gmd\:eastBoundLongitude = "NULL" ;
          		:gmd\:northBoundLatitude = "NULL" ;
          		:gmd\:southBoundLatitude = "NULL" ;
          		:gmd\:westBoundLongitude = "NULL" ;
          		:objectType = "gmd:EX_GeographicBoundingBox" ;
          } // group gmd\:geographicElement
        } // group gmd\:extent

      group: gmd\:characterSet {

        // group attributes:
        		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#MD_CharacterSetCode" ;
        		:codeListValue = "utf8" ;
        		:objectType = "gmd:MD_CharacterSetCode" ;
        } // group gmd\:characterSet

      group: gmd\:descriptiveKeywords {

        // group attributes:
        		:gmd\:keyword = "Atmospheric conditions" ;
        		:objectType = "gmd:MD_Keywords" ;

        group: gmd\:thesaurusName {

          // group attributes:
          		:gmd\:title = "GEMET - INSPIRE themes, version 1.0" ;
          		:objectType = "gmd:CI_Citation" ;

          group: gmd\:date {

            // group attributes:
            		:gmd\:date = "2008-06-01" ;
            		:objectType = "gmd:CI_Date" ;

            group: gmd\:dateType {

              // group attributes:
              		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
              		:codeListValue = "publication" ;
              		:objectType = "gmd:CI_DateTypeCode" ;
              } // group gmd\:dateType
            } // group gmd\:date
          } // group gmd\:thesaurusName

        group: gmd\:type {

          // group attributes:
          		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#MD_KeywordTypeCode" ;
          		:codeListValue = "theme" ;
          		:objectType = "gmd:MD_KeywordTypeCode" ;
          } // group gmd\:type
        } // group gmd\:descriptiveKeywords

      group: gmd\:spatialRepresentationType {

        // group attributes:
        		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#MD_SpatialRepresentationTypeCode" ;
        		:codeListValue = "grid" ;
        		:objectType = "gmd:MD_SpatialRepresentationTypeCode" ;
        } // group gmd\:spatialRepresentationType

      group: gmd\:pointOfContact {

        // group attributes:
        		:gmd\:individualName = "eoHelp" ;
        		:gmd\:organisationName = "Copernicus Space Component Data Access System, ESA, Services Coordinated Interface" ;
        		:gmd\:positionName = "Order Desk" ;
        		:objectType = "gmd:CI_ResponsibleParty" ;

        group: gmd\:contactInfo {

          // group attributes:
          		:objectType = "gmd:CI_Contact" ;

          group: gmd\:address {

            // group attributes:
            		:gmd\:electronicMailAddress = "EOSupport@copernicus.esa.int" ;
            		:objectType = "gmd:CI_Address" ;
            } // group gmd\:address
          } // group gmd\:contactInfo

        group: gmd\:role {

          // group attributes:
          		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_RoleCode" ;
          		:codeListValue = "distributor" ;
          		:objectType = "gmd:CI_RoleCode" ;
          } // group gmd\:role
        } // group gmd\:pointOfContact

      group: gmd\:spatialResolution {

        // group attributes:
        		:gmd\:distance = "7.0" ;
        		:objectType = "gmd:MD_Resolution" ;
        		:uom = "km" ;
        } // group gmd\:spatialResolution
      } // group gmd\:identificationInfo

    group: gmd\:characterSet {

      // group attributes:
      		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#MD_CharacterSetCode" ;
      		:codeListValue = "utf8" ;
      		:objectType = "gmd:MD_CharacterSetCode" ;
      } // group gmd\:characterSet

    group: gmd\:contact {

      // group attributes:
      		:gmd\:individualName = "KNMI Help" ;
      		:gmd\:organisationName = "KNMI" ;
      		:gmd\:positionName = "Help Desk" ;
      		:objectType = "gmd:CI_ResponsibleParty" ;

      group: gmd\:contactInfo {

        // group attributes:
        		:objectType = "gmd:CI_Contact" ;

        group: gmd\:onlineResource {

          // group attributes:
          		:gmd\:function = "information" ;
          		:gmd\:linkage = "http://www.knmi.nl" ;
          		:gmd\:name = "KNMI Home Page" ;
          } // group gmd\:onlineResource

        group: gmd\:address {

          // group attributes:
          		:gmd\:electronicMailAddress = "EOSupport@copernicus.esa.int" ;
          		:objectType = "gmd:CI_Address" ;
          } // group gmd\:address
        } // group gmd\:contactInfo

      group: gmd\:role {

        // group attributes:
        		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_RoleCode" ;
        		:codeListValue = "pointOfContact" ;
        		:objectType = "gmd:CI_RoleCode" ;
        } // group gmd\:role
      } // group gmd\:contact

    group: gmd\:dataQualityInfo {

      // group attributes:
      		:objectType = "gmd:DQ_DataQuality" ;

      group: gmd\:report {

        // group attributes:
        		:objectType = "gmd:DQ_DomainConsistency" ;

        group: gmd\:result {

          // group attributes:
          		:gmd\:pass = "true" ;
          		:gmd\:explanation = "INSPIRE Data specification for orthoimagery is not yet officially published so conformity has not yet been evaluated." ;
          		:objectType = "gmd:DQ_ConformanceResult" ;

          group: gmd\:specification {

            // group attributes:
            		:gmd\:title = "INSPIRE Data Specification on Orthoimagery - Guidelines, version 3.0rc3" ;
            		:objectType = "gmd:CI_Citation" ;

            group: gmd\:date {

              // group attributes:
              		:gmd\:date = "2013-02-04" ;
              		:objectType = "gmd:CI_Date" ;

              group: gmd\:dateType {

                // group attributes:
                		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                		:codeListValue = "publication" ;
                		:objectType = "gmd:CI_DateTypeCode" ;
                } // group gmd\:dateType
              } // group gmd\:date
            } // group gmd\:specification
          } // group gmd\:result
        } // group gmd\:report

      group: gmd\:scope {

        // group attributes:
        		:objectType = "gmd:DQ_Scope" ;

        group: gmd\:level {

          // group attributes:
          		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#MD_ScopeCode" ;
          		:codeListValue = "dataset" ;
          		:objectType = "gmd:MD_ScopeCode" ;
          } // group gmd\:level
        } // group gmd\:scope

      group: gmd\:lineage {

        // group attributes:
        		:objectType = "gmd:LI_Lineage" ;
        		:gmd\:statement = "L1b  dataset produced by the DLR PDGS from the S5p TROPOMI L0 product" ;

        group: gmd\:processStep {

          // group attributes:
          		:gmd\:description = "Processing of L0 to L1b data using the KNMI TROPOMI L01b processor" ;
          		:objectType = "gmi:LE_ProcessStep" ;

          group: gmd\:source\#09 {

            // group attributes:
            		:gmd\:description = "L0 Band 5 NIR science data" ;
            		:objectType = "gmi:LE_Source" ;

            group: gmi\:processedLevel {

              // group attributes:
              		:gmd\:code = "L0" ;
              		:objectType = "gmd:MD_Identifier" ;
              } // group gmi\:processedLevel

            group: gmd\:sourceCitation {

              // group attributes:
              		:objectType = "gmd:CI_Citation" ;

              group: gmd\:date {

                // group attributes:
                		:gmd\:date = "2015-11-18" ;
                		:objectType = "gmd:CI_Date" ;

                group: gmd\:dateType {

                  // group attributes:
                  		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                  		:codeListValue = "creation" ;
                  		:objectType = "gmd:CI_DateTypeCode" ;
                  } // group gmd\:dateType
                } // group gmd\:date

              group: gmd\:title {

                // group attributes:
                		:gco\:characterString = "L0 instrument data for band 5" ;
                } // group gmd\:title

              group: gmd\:alternateTitle\#1 {

                // group attributes:
                		:gmx\:FileName = "S5P_TEST_L0__ODB_4__20140827T114000_20140827T114500_53811_00.RAW" ;
                } // group gmd\:alternateTitle\#1

              group: gmd\:alternateTitle\#2 {

                // group attributes:
                		:gmx\:FileName = "S5P_TEST_L0__ODB_4__20140827T114500_20140827T115000_53811_01.RAW" ;
                } // group gmd\:alternateTitle\#2

              group: gmd\:alternateTitle\#3 {

                // group attributes:
                		:gmx\:FileName = "S5P_TEST_L0__ODB_4__20140827T115000_20140827T115500_53811_02.RAW" ;
                } // group gmd\:alternateTitle\#3

              group: gmd\:alternateTitle\#4 {

                // group attributes:
                		:gmx\:FileName = "S5P_TEST_L0__ODB_4__20140827T115500_20140827T120000_53811_03.RAW" ;
                } // group gmd\:alternateTitle\#4
              } // group gmd\:sourceCitation
            } // group gmd\:source\#09

          group: gmd\:source\#08 {

            // group attributes:
            		:gmd\:description = "L0 Band 4 VIS science data" ;
            		:objectType = "gmi:LE_Source" ;

            group: gmi\:processedLevel {

              // group attributes:
              		:gmd\:code = "L0" ;
              		:objectType = "gmd:MD_Identifier" ;
              } // group gmi\:processedLevel

            group: gmd\:sourceCitation {

              // group attributes:
              		:objectType = "gmd:CI_Citation" ;

              group: gmd\:date {

                // group attributes:
                		:gmd\:date = "2015-11-18" ;
                		:objectType = "gmd:CI_Date" ;

                group: gmd\:dateType {

                  // group attributes:
                  		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                  		:codeListValue = "creation" ;
                  		:objectType = "gmd:CI_DateTypeCode" ;
                  } // group gmd\:dateType
                } // group gmd\:date

              group: gmd\:title {

                // group attributes:
                		:gco\:characterString = "L0 instrument data for band 4" ;
                } // group gmd\:title

              group: gmd\:alternateTitle\#1 {

                // group attributes:
                		:gmx\:FileName = "S5P_TEST_L0__ODB_3__20140827T114000_20140827T114500_53811_00.RAW" ;
                } // group gmd\:alternateTitle\#1

              group: gmd\:alternateTitle\#2 {

                // group attributes:
                		:gmx\:FileName = "S5P_TEST_L0__ODB_3__20140827T114500_20140827T115000_53811_01.RAW" ;
                } // group gmd\:alternateTitle\#2

              group: gmd\:alternateTitle\#3 {

                // group attributes:
                		:gmx\:FileName = "S5P_TEST_L0__ODB_3__20140827T115000_20140827T115500_53811_02.RAW" ;
                } // group gmd\:alternateTitle\#3

              group: gmd\:alternateTitle\#4 {

                // group attributes:
                		:gmx\:FileName = "S5P_TEST_L0__ODB_3__20140827T115500_20140827T120000_53811_03.RAW" ;
                } // group gmd\:alternateTitle\#4
              } // group gmd\:sourceCitation
            } // group gmd\:source\#08

          group: gmd\:source\#11 {

            // group attributes:
            		:gmd\:description = "L0 Band 7 SWIR science data" ;
            		:objectType = "gmi:LE_Source" ;

            group: gmi\:processedLevel {

              // group attributes:
              		:gmd\:code = "L0" ;
              		:objectType = "gmd:MD_Identifier" ;
              } // group gmi\:processedLevel

            group: gmd\:sourceCitation {

              // group attributes:
              		:objectType = "gmd:CI_Citation" ;

              group: gmd\:date {

                // group attributes:
                		:gmd\:date = "2015-11-18" ;
                		:objectType = "gmd:CI_Date" ;

                group: gmd\:dateType {

                  // group attributes:
                  		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                  		:codeListValue = "creation" ;
                  		:objectType = "gmd:CI_DateTypeCode" ;
                  } // group gmd\:dateType
                } // group gmd\:date

              group: gmd\:title {

                // group attributes:
                		:gco\:characterString = "L0 instrument data for band 7" ;
                } // group gmd\:title

              group: gmd\:alternateTitle\#1 {

                // group attributes:
                		:gmx\:FileName = "S5P_TEST_L0__ODB_6__20140827T114000_20140827T114500_53811_00.RAW" ;
                } // group gmd\:alternateTitle\#1

              group: gmd\:alternateTitle\#2 {

                // group attributes:
                		:gmx\:FileName = "S5P_TEST_L0__ODB_6__20140827T114500_20140827T115000_53811_01.RAW" ;
                } // group gmd\:alternateTitle\#2

              group: gmd\:alternateTitle\#3 {

                // group attributes:
                		:gmx\:FileName = "S5P_TEST_L0__ODB_6__20140827T115000_20140827T115500_53811_02.RAW" ;
                } // group gmd\:alternateTitle\#3

              group: gmd\:alternateTitle\#4 {

                // group attributes:
                		:gmx\:FileName = "S5P_TEST_L0__ODB_6__20140827T115500_20140827T120000_53811_03.RAW" ;
                } // group gmd\:alternateTitle\#4
              } // group gmd\:sourceCitation
            } // group gmd\:source\#11

          group: gmd\:source\#01 {

            // group attributes:
            		:gmd\:description = "Auxiliary Calibration Key Data product" ;
            		:objectType = "gmi:LE_Source" ;

            group: gmd\:sourceCitation {

              // group attributes:
              		:objectType = "gmd:CI_Citation" ;

              group: gmd\:date {

                // group attributes:
                		:gmd\:date = "2015-11-18" ;
                		:objectType = "gmd:CI_Date" ;

                group: gmd\:dateType {

                  // group attributes:
                  		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                  		:codeListValue = "creation" ;
                  		:objectType = "gmd:CI_DateTypeCode" ;
                  } // group gmd\:dateType
                } // group gmd\:date

              group: gmd\:title {

                // group attributes:
                		:gco\:characterString = "Auxiliary Calibration Key Data Set" ;
                } // group gmd\:title

              group: gmd\:alternateTitle\#1 {

                // group attributes:
                		:gmx\:FileName = "S5P_TEST_AUX_L1_CKD_20140101T000000_20151231T000000_00000_01_000900_20150915T120000.h5" ;
                } // group gmd\:alternateTitle\#1
              } // group gmd\:sourceCitation
            } // group gmd\:source\#01

          group: gmd\:source\#13 {

            // group attributes:
            		:gmd\:description = "L0 Ancillary data" ;
            		:objectType = "gmi:LE_Source" ;

            group: gmi\:processedLevel {

              // group attributes:
              		:gmd\:code = "L0" ;
              		:objectType = "gmd:MD_Identifier" ;
              } // group gmi\:processedLevel

            group: gmd\:sourceCitation {

              // group attributes:
              		:objectType = "gmd:CI_Citation" ;

              group: gmd\:date {

                // group attributes:
                		:gmd\:date = "2015-11-18" ;
                		:objectType = "gmd:CI_Date" ;

                group: gmd\:dateType {

                  // group attributes:
                  		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                  		:codeListValue = "creation" ;
                  		:objectType = "gmd:CI_DateTypeCode" ;
                  } // group gmd\:dateType
                } // group gmd\:date

              group: gmd\:title {

                // group attributes:
                		:gco\:characterString = "L0 instrument ancillary data" ;
                } // group gmd\:title

              group: gmd\:alternateTitle\#1 {

                // group attributes:
                		:gmx\:FileName = "S5P_TEST_L0__SAT_A__20140827T114000_20140827T114500_53811_00.RAW" ;
                } // group gmd\:alternateTitle\#1

              group: gmd\:alternateTitle\#2 {

                // group attributes:
                		:gmx\:FileName = "S5P_TEST_L0__SAT_A__20140827T114500_20140827T115000_53811_01.RAW" ;
                } // group gmd\:alternateTitle\#2

              group: gmd\:alternateTitle\#3 {

                // group attributes:
                		:gmx\:FileName = "S5P_TEST_L0__SAT_A__20140827T115000_20140827T115500_53811_02.RAW" ;
                } // group gmd\:alternateTitle\#3

              group: gmd\:alternateTitle\#4 {

                // group attributes:
                		:gmx\:FileName = "S5P_TEST_L0__SAT_A__20140827T115500_20140827T120000_53811_03.RAW" ;
                } // group gmd\:alternateTitle\#4
              } // group gmd\:sourceCitation
            } // group gmd\:source\#13

          group: gmd\:source\#03 {

            group: gmd\:sourceCitation {

              // group attributes:
              		:objectType = "gmd:CI_Citation" ;

              group: gmd\:date {

                // group attributes:
                		:gmd\:date = "2015-11-18" ;
                		:objectType = "gmd:CI_Date" ;

                group: gmd\:dateType {

                  // group attributes:
                  		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                  		:codeListValue = "creation" ;
                  		:objectType = "gmd:CI_DateTypeCode" ;
                  } // group gmd\:dateType
                } // group gmd\:date

              group: gmd\:title {

                // group attributes:
                		:gco\:characterString = "In-flight Calibration Key Data Set UVN" ;
                } // group gmd\:title

              group: gmd\:alternateTitle\#1 {

                // group attributes:
                		:gmx\:FileName = "S5P_TEST_ICM_CKDSIR_20140101T000000_20151231T000000_00000_01_000900_20150915T120000.h5" ;
                } // group gmd\:alternateTitle\#1
              } // group gmd\:sourceCitation
            } // group gmd\:source\#03

          group: gmd\:source\#02 {

            // group attributes:
            		:gmd\:description = "In-flight UVN Calibration Key Data product" ;
            		:objectType = "gmi:LE_Source" ;

            group: gmd\:sourceCitation {

              // group attributes:
              		:objectType = "gmd:CI_Citation" ;

              group: gmd\:date {

                // group attributes:
                		:gmd\:date = "2015-11-18" ;
                		:objectType = "gmd:CI_Date" ;

                group: gmd\:dateType {

                  // group attributes:
                  		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                  		:codeListValue = "creation" ;
                  		:objectType = "gmd:CI_DateTypeCode" ;
                  } // group gmd\:dateType
                } // group gmd\:date

              group: gmd\:title {

                // group attributes:
                		:gco\:characterString = "In-flight Calibration Key Data Set UVN" ;
                } // group gmd\:title

              group: gmd\:alternateTitle\#1 {

                // group attributes:
                		:gmx\:FileName = "S5P_TEST_ICM_CKDUVN_20140101T000000_20151231T000000_00000_01_000900_20150915T120000.h5" ;
                } // group gmd\:alternateTitle\#1
              } // group gmd\:sourceCitation
            } // group gmd\:source\#02

          group: gmd\:source\#05 {

            // group attributes:
            		:gmd\:description = "L0 Band 1 UV science data" ;
            		:objectType = "gmi:LE_Source" ;

            group: gmi\:processedLevel {

              // group attributes:
              		:gmd\:code = "L0" ;
              		:objectType = "gmd:MD_Identifier" ;
              } // group gmi\:processedLevel

            group: gmd\:sourceCitation {

              // group attributes:
              		:objectType = "gmd:CI_Citation" ;

              group: gmd\:date {

                // group attributes:
                		:gmd\:date = "2015-11-18" ;
                		:objectType = "gmd:CI_Date" ;

                group: gmd\:dateType {

                  // group attributes:
                  		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                  		:codeListValue = "creation" ;
                  		:objectType = "gmd:CI_DateTypeCode" ;
                  } // group gmd\:dateType
                } // group gmd\:date

              group: gmd\:title {

                // group attributes:
                		:gco\:characterString = "L0 instrument data for band 1" ;
                } // group gmd\:title

              group: gmd\:alternateTitle\#1 {

                // group attributes:
                		:gmx\:FileName = "S5P_TEST_L0__ODB_8__20140827T114000_20140827T114500_53811_00.RAW" ;
                } // group gmd\:alternateTitle\#1

              group: gmd\:alternateTitle\#2 {

                // group attributes:
                		:gmx\:FileName = "S5P_TEST_L0__ODB_8__20140827T114500_20140827T115000_53811_01.RAW" ;
                } // group gmd\:alternateTitle\#2

              group: gmd\:alternateTitle\#3 {

                // group attributes:
                		:gmx\:FileName = "S5P_TEST_L0__ODB_8__20140827T115000_20140827T115500_53811_02.RAW" ;
                } // group gmd\:alternateTitle\#3

              group: gmd\:alternateTitle\#4 {

                // group attributes:
                		:gmx\:FileName = "S5P_TEST_L0__ODB_8__20140827T115500_20140827T120000_53811_03.RAW" ;
                } // group gmd\:alternateTitle\#4
              } // group gmd\:sourceCitation
            } // group gmd\:source\#05

          group: gmd\:source\#04 {

            // group attributes:
            		:gmd\:description = "L0 Engineering data" ;
            		:objectType = "gmi:LE_Source" ;

            group: gmi\:processedLevel {

              // group attributes:
              		:gmd\:code = "L0" ;
              		:objectType = "gmd:MD_Identifier" ;
              } // group gmi\:processedLevel

            group: gmd\:sourceCitation {

              // group attributes:
              		:objectType = "gmd:CI_Citation" ;

              group: gmd\:date {

                // group attributes:
                		:gmd\:date = "2015-11-18" ;
                		:objectType = "gmd:CI_Date" ;

                group: gmd\:dateType {

                  // group attributes:
                  		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                  		:codeListValue = "creation" ;
                  		:objectType = "gmd:CI_DateTypeCode" ;
                  } // group gmd\:dateType
                } // group gmd\:date

              group: gmd\:title {

                // group attributes:
                		:gco\:characterString = "L0 instrument engineering data" ;
                } // group gmd\:title

              group: gmd\:alternateTitle\#1 {

                // group attributes:
                		:gmx\:FileName = "S5P_TEST_L0__ENG_A__20140827T114000_20140827T114500_53811_00.RAW" ;
                } // group gmd\:alternateTitle\#1

              group: gmd\:alternateTitle\#2 {

                // group attributes:
                		:gmx\:FileName = "S5P_TEST_L0__ENG_A__20140827T114500_20140827T115000_53811_01.RAW" ;
                } // group gmd\:alternateTitle\#2

              group: gmd\:alternateTitle\#3 {

                // group attributes:
                		:gmx\:FileName = "S5P_TEST_L0__ENG_A__20140827T115000_20140827T115500_53811_02.RAW" ;
                } // group gmd\:alternateTitle\#3

              group: gmd\:alternateTitle\#4 {

                // group attributes:
                		:gmx\:FileName = "S5P_TEST_L0__ENG_A__20140827T115500_20140827T120000_53811_03.RAW" ;
                } // group gmd\:alternateTitle\#4
              } // group gmd\:sourceCitation
            } // group gmd\:source\#04

          group: gmd\:source\#07 {

            // group attributes:
            		:gmd\:description = "L0 Band 3 VIS science data" ;
            		:objectType = "gmi:LE_Source" ;

            group: gmi\:processedLevel {

              // group attributes:
              		:gmd\:code = "L0" ;
              		:objectType = "gmd:MD_Identifier" ;
              } // group gmi\:processedLevel

            group: gmd\:sourceCitation {

              // group attributes:
              		:objectType = "gmd:CI_Citation" ;

              group: gmd\:date {

                // group attributes:
                		:gmd\:date = "2015-11-18" ;
                		:objectType = "gmd:CI_Date" ;

                group: gmd\:dateType {

                  // group attributes:
                  		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                  		:codeListValue = "creation" ;
                  		:objectType = "gmd:CI_DateTypeCode" ;
                  } // group gmd\:dateType
                } // group gmd\:date

              group: gmd\:title {

                // group attributes:
                		:gco\:characterString = "L0 instrument data for band 3" ;
                } // group gmd\:title

              group: gmd\:alternateTitle\#1 {

                // group attributes:
                		:gmx\:FileName = "S5P_TEST_L0__ODB_2__20140827T114000_20140827T114500_53811_00.RAW" ;
                } // group gmd\:alternateTitle\#1

              group: gmd\:alternateTitle\#2 {

                // group attributes:
                		:gmx\:FileName = "S5P_TEST_L0__ODB_2__20140827T114500_20140827T115000_53811_01.RAW" ;
                } // group gmd\:alternateTitle\#2

              group: gmd\:alternateTitle\#3 {

                // group attributes:
                		:gmx\:FileName = "S5P_TEST_L0__ODB_2__20140827T115000_20140827T115500_53811_02.RAW" ;
                } // group gmd\:alternateTitle\#3

              group: gmd\:alternateTitle\#4 {

                // group attributes:
                		:gmx\:FileName = "S5P_TEST_L0__ODB_2__20140827T115500_20140827T120000_53811_03.RAW" ;
                } // group gmd\:alternateTitle\#4
              } // group gmd\:sourceCitation
            } // group gmd\:source\#07

          group: gmd\:source\#06 {

            // group attributes:
            		:gmd\:description = "L0 Band 2 UV science data" ;
            		:objectType = "gmi:LE_Source" ;

            group: gmi\:processedLevel {

              // group attributes:
              		:gmd\:code = "L0" ;
              		:objectType = "gmd:MD_Identifier" ;
              } // group gmi\:processedLevel

            group: gmd\:sourceCitation {

              // group attributes:
              		:objectType = "gmd:CI_Citation" ;

              group: gmd\:date {

                // group attributes:
                		:gmd\:date = "2015-11-18" ;
                		:objectType = "gmd:CI_Date" ;

                group: gmd\:dateType {

                  // group attributes:
                  		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                  		:codeListValue = "creation" ;
                  		:objectType = "gmd:CI_DateTypeCode" ;
                  } // group gmd\:dateType
                } // group gmd\:date

              group: gmd\:title {

                // group attributes:
                		:gco\:characterString = "L0 instrument data for band 2" ;
                } // group gmd\:title

              group: gmd\:alternateTitle\#1 {

                // group attributes:
                		:gmx\:FileName = "S5P_TEST_L0__ODB_1__20140827T114000_20140827T114500_53811_00.RAW" ;
                } // group gmd\:alternateTitle\#1

              group: gmd\:alternateTitle\#2 {

                // group attributes:
                		:gmx\:FileName = "S5P_TEST_L0__ODB_1__20140827T114500_20140827T115000_53811_01.RAW" ;
                } // group gmd\:alternateTitle\#2

              group: gmd\:alternateTitle\#3 {

                // group attributes:
                		:gmx\:FileName = "S5P_TEST_L0__ODB_1__20140827T115000_20140827T115500_53811_02.RAW" ;
                } // group gmd\:alternateTitle\#3

              group: gmd\:alternateTitle\#4 {

                // group attributes:
                		:gmx\:FileName = "S5P_TEST_L0__ODB_1__20140827T115500_20140827T120000_53811_03.RAW" ;
                } // group gmd\:alternateTitle\#4
              } // group gmd\:sourceCitation
            } // group gmd\:source\#06

          group: gmd\:source\#12 {

            // group attributes:
            		:gmd\:description = "L0 Band 8 SWIR science data" ;
            		:objectType = "gmi:LE_Source" ;

            group: gmi\:processedLevel {

              // group attributes:
              		:gmd\:code = "L0" ;
              		:objectType = "gmd:MD_Identifier" ;
              } // group gmi\:processedLevel

            group: gmd\:sourceCitation {

              // group attributes:
              		:objectType = "gmd:CI_Citation" ;

              group: gmd\:date {

                // group attributes:
                		:gmd\:date = "2015-11-18" ;
                		:objectType = "gmd:CI_Date" ;

                group: gmd\:dateType {

                  // group attributes:
                  		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                  		:codeListValue = "creation" ;
                  		:objectType = "gmd:CI_DateTypeCode" ;
                  } // group gmd\:dateType
                } // group gmd\:date

              group: gmd\:title {

                // group attributes:
                		:gco\:characterString = "L0 instrument data for band 8" ;
                } // group gmd\:title

              group: gmd\:alternateTitle\#1 {

                // group attributes:
                		:gmx\:FileName = "S5P_TEST_L0__ODB_7__20140827T114000_20140827T114500_53811_00.RAW" ;
                } // group gmd\:alternateTitle\#1

              group: gmd\:alternateTitle\#2 {

                // group attributes:
                		:gmx\:FileName = "S5P_TEST_L0__ODB_7__20140827T114500_20140827T115000_53811_01.RAW" ;
                } // group gmd\:alternateTitle\#2

              group: gmd\:alternateTitle\#3 {

                // group attributes:
                		:gmx\:FileName = "S5P_TEST_L0__ODB_7__20140827T115000_20140827T115500_53811_02.RAW" ;
                } // group gmd\:alternateTitle\#3

              group: gmd\:alternateTitle\#4 {

                // group attributes:
                		:gmx\:FileName = "S5P_TEST_L0__ODB_7__20140827T115500_20140827T120000_53811_03.RAW" ;
                } // group gmd\:alternateTitle\#4
              } // group gmd\:sourceCitation
            } // group gmd\:source\#12

          group: gmi\:report {

            // group attributes:
            		:gmi\:description = "L0 processed to L1b data using the KNMI TROPOMI L01b processor" ;
            		:gmi\:fileType = "netCDF" ;
            		:gmi\:name = "TROPOMI L01b processing report" ;
            		:objectType = "gmi:LE_ProcessStepReport" ;
            } // group gmi\:report

          group: gmi\:processingInformation {

            // group attributes:
            		:objectType = "gmi:LE_Processing" ;

            group: gmi\:softwareReference {

              // group attributes:
              		:gmd\:title = "L01b processor description" ;
              		:objectType = "gmd:CI_Citation" ;

              group: gmd\:date {

                // group attributes:
                		:gmd\:date = "2014-12-31" ;
                		:objectType = "gmd:CI_Date" ;

                group: gmd\:dateType {

                  // group attributes:
                  		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                  		:codeListValue = "creation" ;
                  		:objectType = "gmd:CI_DateTypeCode" ;
                  } // group gmd\:dateType
                } // group gmd\:date
              } // group gmi\:softwareReference

            group: gmi\:documentation\#1 {

              // group attributes:
              		:objectType = "gmd:CI_Citation" ;
              		:gmd\:title = "S5P-KNMI-L01B-0009-SD-algorithm_theoretical_basis_document-3.0.0-20140707.pdf" ;

              group: gmd\:date {

                // group attributes:
                		:gmd\:date = "2014-07-07" ;
                		:objectType = "gmd:CI_Date" ;

                group: gmd\:dateType {

                  // group attributes:
                  		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                  		:codeListValue = "publication" ;
                  		:objectType = "gmd:CI_DateTypeCode" ;
                  } // group gmd\:dateType
                } // group gmd\:date
              } // group gmi\:documentation\#1

            group: gmi\:identifier {

              // group attributes:
              		:gmd\:code = "KNMI TROPOMI L01b processor" ;
              		:objectType = "gmd:MD_Identifier" ;
              } // group gmi\:identifier

            group: gmi\:documentation\#2 {

              // group attributes:
              		:gmd\:title = "S5P-KNMI-L01B-0012-SD-input_output_data_specification-3.0.0-20140707.pdf" ;
              		:objectType = "gmd:CI_Citation" ;

              group: gmd\:date {

                // group attributes:
                		:gmd\:date = "2014-07-07" ;
                		:objectType = "gmd:CI_Date" ;

                group: gmd\:dateType {

                  // group attributes:
                  		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                  		:codeListValue = "publication" ;
                  		:objectType = "gmd:CI_DateTypeCode" ;
                  } // group gmd\:dateType
                } // group gmd\:date
              } // group gmi\:documentation\#2
            } // group gmi\:processingInformation

          group: gmi\:output {

            // group attributes:
            		:gmd\:description = "TROPOMI L1b Radiance product band 6 (NIR detector)" ;
            		:objectType = "gmi:LE_Source" ;

            group: gmi\:processedLevel {

              // group attributes:
              		:gmd\:code = "L1b" ;
              		:objectType = "gmd:MD_Identifier" ;
              } // group gmi\:processedLevel

            group: gmd\:sourceCitation {

              // group attributes:
              		:objectType = "gmd:CI_Citation" ;
              		:gmd\:title = "S5P_TEST_L1B_RA_BD6_20140827T114200_20140827T115800_53811_01_000901_20141209T120000" ;

              group: gmd\:date {

                // group attributes:
                		:gmd\:date = "2015-11-18" ;
                		:objectType = "gmd:CI_Date" ;

                group: gmd\:dateType {

                  // group attributes:
                  		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                  		:codeListValue = "creation" ;
                  		:objectType = "gmd:CI_DateTypeCode" ;
                  } // group gmd\:dateType
                } // group gmd\:date
              } // group gmd\:sourceCitation
            } // group gmi\:output

          group: gmd\:source\#10 {

            // group attributes:
            		:gmd\:description = "L0 Band 6 NIR science data" ;
            		:objectType = "gmi:LE_Source" ;

            group: gmi\:processedLevel {

              // group attributes:
              		:gmd\:code = "L0" ;
              		:objectType = "gmd:MD_Identifier" ;
              } // group gmi\:processedLevel

            group: gmd\:sourceCitation {

              // group attributes:
              		:objectType = "gmd:CI_Citation" ;

              group: gmd\:date {

                // group attributes:
                		:gmd\:date = "2015-11-18" ;
                		:objectType = "gmd:CI_Date" ;

                group: gmd\:dateType {

                  // group attributes:
                  		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                  		:codeListValue = "creation" ;
                  		:objectType = "gmd:CI_DateTypeCode" ;
                  } // group gmd\:dateType
                } // group gmd\:date

              group: gmd\:title {

                // group attributes:
                		:gco\:characterString = "L0 instrument data for band 6" ;
                } // group gmd\:title

              group: gmd\:alternateTitle\#1 {

                // group attributes:
                		:gmx\:FileName = "S5P_TEST_L0__ODB_5__20140827T114000_20140827T114500_53811_00.RAW" ;
                } // group gmd\:alternateTitle\#1

              group: gmd\:alternateTitle\#2 {

                // group attributes:
                		:gmx\:FileName = "S5P_TEST_L0__ODB_5__20140827T114500_20140827T115000_53811_01.RAW" ;
                } // group gmd\:alternateTitle\#2

              group: gmd\:alternateTitle\#3 {

                // group attributes:
                		:gmx\:FileName = "S5P_TEST_L0__ODB_5__20140827T115000_20140827T115500_53811_02.RAW" ;
                } // group gmd\:alternateTitle\#3

              group: gmd\:alternateTitle\#4 {

                // group attributes:
                		:gmx\:FileName = "S5P_TEST_L0__ODB_5__20140827T115500_20140827T120000_53811_03.RAW" ;
                } // group gmd\:alternateTitle\#4
              } // group gmd\:sourceCitation
            } // group gmd\:source\#10
          } // group gmd\:processStep
        } // group gmd\:lineage
      } // group gmd\:dataQualityInfo

    group: gmd\:language {

      // group attributes:
      		:codeList = "http://www.loc.gov/standards/iso639-2/" ;
      		:codeListValue = "eng" ;
      		:objectType = "gmd:LanguageCode" ;
      } // group gmd\:language
    } // group ISO_METADATA
  } // group METADATA

group: PROCESSOR {
  dimensions:
  	algorithm_configuration_dim = 313 ;
  	job_configuration_dim = 136 ;
  	processing_configuration_dim = 1410 ;
  variables:
  	string algorithm_configuration(algorithm_configuration_dim) ;
  		algorithm_configuration:description = "Overview of the algorithms that were used in de L01b data processing for this data product" ;
  	string job_configuration(job_configuration_dim) ;
  		job_configuration:description = "Internal representation of the job configuration of the L01b data processing for this data product" ;
  	string processing_configuration(processing_configuration_dim) ;
  		processing_configuration:description = "Overview of all the processing steps, the algorithm order and data flow of the L01b data processing for this data product" ;
  } // group PROCESSOR
}
