netcdf car-dim {
dimensions:
	time = 22951 ;
	NumberOfChannels = 14 ;
	angel = 361 ;
variables:
	int Date(time) ;
		Date:long_name = "Date" ;
		Date:Data_Aquistion_Date = "YYYYMMDD" ;
		Date:origname = "Date" ;
		Date:_ChunkSizes = 22951 ;
	float CoordinatedUniversalTime(time) ;
		CoordinatedUniversalTime:UTC_time = "HHMMSS.S" ;
		CoordinatedUniversalTime:origname = "CoordinatedUniversalTime" ;
		CoordinatedUniversalTime:long_name = "CoordinatedUniversalTime" ;
		CoordinatedUniversalTime:_ChunkSizes = 22951 ;
	float GPSAltitude(time) ;
		GPSAltitude:GPS_height = "GPS height Meter " ;
		GPSAltitude:origname = "GPSAltitude" ;
		GPSAltitude:long_name = "GPSAltitude" ;
		GPSAltitude:_ChunkSizes = 22951 ;
	float AircraftLatitude(time) ;
		AircraftLatitude:Latitude = "Aircraft Latitude Degrees" ;
		AircraftLatitude:origname = "AircraftLatitude" ;
		AircraftLatitude:long_name = "AircraftLatitude" ;
		AircraftLatitude:_ChunkSizes = 22951 ;
	float AircraftLongitude(time) ;
		AircraftLongitude:Longitude = "Aircraft Longitude Degrees" ;
		AircraftLongitude:origname = "AircraftLongitude" ;
		AircraftLongitude:long_name = "AircraftLongitude" ;
		AircraftLongitude:_ChunkSizes = 22951 ;
	float AircraftHeading(time) ;
		AircraftHeading:long_name = "AircraftHeading" ;
		AircraftHeading:Heading = "Aircraft Heading Degrees" ;
		AircraftHeading:origname = "AircraftHeading" ;
		AircraftHeading:_ChunkSizes = 22951 ;
	float AircraftPitch(time) ;
		AircraftPitch:Aircraft_Pitch = "Aircraft Pitch Degrees " ;
		AircraftPitch:origname = "AircraftPitch" ;
		AircraftPitch:long_name = "AircraftPitch" ;
		AircraftPitch:_ChunkSizes = 22951 ;
	int ScanLineCounter(time) ;
		ScanLineCounter:scan_line_count = "Scan lines from data start" ;
		ScanLineCounter:origname = "ScanLineCounter" ;
		ScanLineCounter:long_name = "ScanLineCounter" ;
		ScanLineCounter:_ChunkSizes = 22951 ;
	double lambda_340nm(time, angel) ;
		lambda_340nm:CAR_ch1 = "0.340 reflectance 0.5 degree interval" ;
		lambda_340nm:origname = "lambda_340nm" ;
		lambda_340nm:long_name = "lambda_340nm" ;
		lambda_340nm:_ChunkSizes = 5738, 73 ;
	double lambda_380nm(time, angel) ;
		lambda_380nm:CAR_ch2 = "0.381 reflectance 0.5 degree interval" ;
		lambda_380nm:origname = "lambda_380nm" ;
		lambda_380nm:long_name = "lambda_380nm" ;
		lambda_380nm:_ChunkSizes = 5738, 73 ;
	double lambda_470nm(time, angel) ;
		lambda_470nm:CAR_ch3 = "0.472 reflectance 0.5 degree interval" ;
		lambda_470nm:origname = "lambda_470nm" ;
		lambda_470nm:long_name = "lambda_470nm" ;
		lambda_470nm:_ChunkSizes = 5738, 73 ;
	double lambda_680nm(time, angel) ;
		lambda_680nm:CAR_ch4 = "0.682 reflectance 0.5 degree interval" ;
		lambda_680nm:origname = "lambda_680nm" ;
		lambda_680nm:long_name = "lambda_680nm" ;
		lambda_680nm:_ChunkSizes = 5738, 73 ;
	double lambda_870nm(time, angel) ;
		lambda_870nm:CAR_ch5 = "0.870 reflectance 0.5 degree interval" ;
		lambda_870nm:origname = "lambda_870nm" ;
		lambda_870nm:long_name = "lambda_870nm" ;
		lambda_870nm:_ChunkSizes = 5738, 73 ;
	double lambda_1037nm(time, angel) ;
		lambda_1037nm:CAR_ch6 = "1.036 reflectance 0.5 degree interval" ;
		lambda_1037nm:origname = "lambda_1037nm" ;
		lambda_1037nm:long_name = "lambda_1037nm" ;
		lambda_1037nm:_ChunkSizes = 5738, 73 ;
	double lambda_610nm(time, angel) ;
		lambda_610nm:CAR_ch7 = "0.610 reflectance 0.5 degree interval" ;
		lambda_610nm:origname = "lambda_610nm" ;
		lambda_610nm:long_name = "lambda_610nm" ;
		lambda_610nm:_ChunkSizes = 5738, 73 ;
	double lambda_1275nm(time, angel) ;
		lambda_1275nm:CAR_ch8 = "1.273 reflectance 0.5 degree interval" ;
		lambda_1275nm:origname = "lambda_1275nm" ;
		lambda_1275nm:long_name = "lambda_1275nm" ;
		lambda_1275nm:_ChunkSizes = 5738, 73 ;
	double lambda_1564nm(time, angel) ;
		lambda_1564nm:CAR_ch9 = "1.562 reflectance 0.5 degree interval" ;
		lambda_1564nm:origname = "lambda_1564nm" ;
		lambda_1564nm:long_name = "lambda_1564nm" ;
		lambda_1564nm:_ChunkSizes = 5738, 73 ;
	double lambda_1657nm(time, angel) ;
		lambda_1657nm:CAR_ch10 = "1.656 reflectance 0.5 degree interval" ;
		lambda_1657nm:origname = "lambda_1657nm" ;
		lambda_1657nm:long_name = "lambda_1657nm" ;
		lambda_1657nm:_ChunkSizes = 5738, 73 ;
	double lambda_1738nm(time, angel) ;
		lambda_1738nm:CAR_ch11 = "1.737 reflectance 0.5 degree interval" ;
		lambda_1738nm:origname = "lambda_1738nm" ;
		lambda_1738nm:long_name = "lambda_1738nm" ;
		lambda_1738nm:_ChunkSizes = 5738, 73 ;
	double lambda_2105nm(time, angel) ;
		lambda_2105nm:CAR_ch12 = "2.103 reflectance 0.5 degree interval" ;
		lambda_2105nm:origname = "lambda_2105nm" ;
		lambda_2105nm:long_name = "lambda_2105nm" ;
		lambda_2105nm:_ChunkSizes = 5738, 73 ;
	double lambda_2202nm(time, angel) ;
		lambda_2202nm:CAR_ch13 = "2.205 reflectance 0.5 degree interval" ;
		lambda_2202nm:origname = "lambda_2202nm" ;
		lambda_2202nm:long_name = "lambda_2202nm" ;
		lambda_2202nm:_ChunkSizes = 5738, 73 ;
	double lambda_2303nm(time, angel) ;
		lambda_2303nm:CAR_ch14 = "2.301 reflectance 0.5 degree interval" ;
		lambda_2303nm:origname = "lambda_2303nm" ;
		lambda_2303nm:long_name = "lambda_2303nm" ;
		lambda_2303nm:_ChunkSizes = 5738, 73 ;
	float SolarZenithAngle(time) ;
		SolarZenithAngle:Solar_Zenith = "Solar Zenith Angle Degrees" ;
		SolarZenithAngle:origname = "SolarZenithAngle" ;
		SolarZenithAngle:long_name = "SolarZenithAngle" ;
		SolarZenithAngle:_ChunkSizes = 22951 ;
	float SolarAzimuthAngle(time) ;
		SolarAzimuthAngle:Solar_Azimuth = "Solar Azimuth Angle Degrees" ;
		SolarAzimuthAngle:origname = "SolarAzimuthAngle" ;
		SolarAzimuthAngle:long_name = "SolarAzimuthAngle" ;
		SolarAzimuthAngle:_ChunkSizes = 22951 ;
	float CentralWavelength(NumberOfChannels) ;
		CentralWavelength:CentralWavelength = "CAR Channel CentralWavelength" ;
		CentralWavelength:origname = "CentralWavelength" ;
		CentralWavelength:long_name = "CentralWavelength" ;
		CentralWavelength:_ChunkSizes = 14 ;
	int SolarIrradiance(NumberOfChannels) ;
		SolarIrradiance:Solar_Spectral_irridiance = "Solar Spectral Irridiance for each channel" ;
		SolarIrradiance:origname = "SolarIrradiance" ;
		SolarIrradiance:long_name = "SolarIrradiance" ;
		SolarIrradiance:_ChunkSizes = 14 ;

// global attributes:
		:Version = "CAR level 1C product" ;
		:Date = "Jun 25,2015" ;
		:Experiment_Name = "Discover AQ" ;
		:Instrument_PI = "Charles K. Gatebe" ;
		:email = "charles.k.gatebe@nasa.gov" ;
		:Website = "http://car.gsfc.nasa.gov" ;
}
