// Contributed by Jessica Hausman <Jessica.K.Hausman AT jpl DOT nasa DOT gov>

netcdf Q2014050173000.L2_SCI_V4 {

// global attributes:
		:Product\ Name = "Q2014050173000.L2_SCI_V4.0" ;
		:Title = "Aquarius Level 2 Data" ;
		:Data\ Center = "NASA/GSFC Aquarius Data Processing Center" ;
		:Mission = "SAC-D Aquarius" ;
		:Mission\ Characteristics = "Nominal orbit: inclination=98.0 (Sun-synchronous); node=6PM (ascending); eccentricity=<0.002; altitude=657 km; ground speed=6.825 km/sec" ;
		:Sensor = "Aquarius" ;
		:Sensor\ Characteristics = "Number of beams=3; channels per receiver=4; frequency 1.413 GHz; bits per sample=16; instatntaneous field of view=6.5 degrees; science data block period=1.44 sec." ;
		:Data\ Type = "SCI" ;
		:Software\ ID = "4.00" ;
		:Processing\ Version = "V4.0" ;
		:Processing\ Time = "2015155172224000" ;
		:Input\ Files = "Q2014050173000.L1A_SCI" ;
		:Processing\ Control = "ifile=/data7/sdpsoper/vdc/vpu6/workbuf/Q2014050173000.L1A_SCI ofile=/data7/sdpsoper/vdc/vpu6/workbuf/Q2014050173000.L2_SCI_V4.0 yancfile1=y2014021912.h5 yancfile2=y2014021918.h5 yancfile3=y2014022000.h5 c_delta_TND=0.005957319097863 0.012382688000750 0.000688525722399 0.005498736477495 0.009869297059855 0.000587055056684 0.006316487443884 0.013593252195015 0.000713618469860 0.005016272510612 0.010186625543718 0.000650544867204 0.006233499611709 0.009903518037236 0.000529897823645 0.006068613199395 0.010888564961881 0.000618946224004 ta_nominal_files=$OCDATAROOT/aquarius/radiometer/Ta_nom_4Apr2014_v2.lst wind_errortab_file=$OCDATAROOT/aquarius/radiometer/error_tab.h5 emiss_coeff_harm_file=$OCDATAROOT/aquarius/radiometer/deW_harm_coeffs_V9A_MI.h5 scat_coeff_harm_file=$OCDATAROOT/aquarius/radiometer/sigma0_harm_coeffs_V9A_MI.h5 climate_sal_file=$OCDATAROOT/aquarius/radiometer/AQ_SSS_clim_map_testbedV41_2year.h5 dtbw_win_sigma_file=$OCDATAROOT/aquarius/radiometer/dtbw_residual_win_sigma_bin_flag_V9_HHH_A.h5 dtbw_win_wav_file=$OCDATAROOT/aquarius/radiometer/dtbw_residual_win_wav_bin_V9_HHH_A.h5 rad_dta_gal_file=$OCDATAROOT/aquarius/radiometer/dta_gal_symm.h5 sss_algorithm=SIGMA0_HHH l2prod=default:rad_hh_wind_speed,rad_hhh_wind_speed,rad_exp_TaV_hhh,rad_exp_TaH_hhh,rad_exp_Ta3_hhh,anc_swh,rad_galact_Ta_ref_GO_V,rad_galact_Ta_ref_GO_H,rad_galact_dTa_V,rad_galact_dTa_H,rad_dtb_sst_wspd_V,rad_dtb_sst_wspd_H,density,SSS_unc_ran,SSS_unc_sys rad_offset_corr_file=$OCVARROOT/aquarius/rad_offset_corr_V400_Liang.h5 rad_apc_file=$OCDATAROOT/aquarius/radiometer/apc_matrix_may2013_1.h5 coeff_loss_file=$OCDATAROOT/aquarius/radiometer/coeff_loss_V4.txt rfi_mask_file=$OCDATAROOT/aquarius/radiometer/rfi_mask_1.h5 radflaglimitsfile=$OCDATAROOT/aquarius/radiometer/radiometer_flag_limits.txt dtb_emiss_wspd_file=$OCDATAROOT/aquarius/radiometer/dtb_emiss_wspd.h5 dI_U_coeff_file=$OCDATAROOT/aquarius/radiometer/dI_U_fit.h5 l2_uncertainty_maps_file=$OCDATAROOT/aquarius/radiometer/L2_uncertainty_maps_AD_V4.0.h5 rad_gainice_file=$OCDATAROOT/aquarius/radiometer/gain_ice_V3.6.h5 rad_landcorr_file=$OCDATAROOT/aquarius/radiometer/land_corr_tables_V3.6.h5 rad_landtables_file=$OCDATAROOT/aquarius/radiometer/land_tables_V3.6.h5 rad_sun_file=$OCDATAROOT/aquarius/radiometer/sun_tables_V3.6.h5 pversion=V4.0 xrayfile1=/data7/sdpsoper/vdc/vpu6/workbuf/N201405000_XRAY_GOES_24h.h5 rad_tausq_file=$OCDATAROOT/aquarius/radiometer/tausq.h5 rad_sunbak_file=$OCDATAROOT/aquarius/radiometer/sun_bak_tables.h5 rad_oceanrefl_file=$OCDATAROOT/aquarius/radiometer/ocean_reflectance.h5 rad_galwind_file=$OCDATAROOT/aquarius/radiometer/galaxy_wind_tables_V2.0.h5 coeff_nl_file=$OCDATAROOT/aquarius/radiometer/coeff_nl.txt matchup_lat=-999 matchup_lon=-999 matchup_delta_lat=1.0 matchup_delta_lon=1.0 matchup_min_distance=35.0 browse=false iopt_rfi=true iopt_nosa1=true iopt_l1b=false matchup_limits_file= rpy_adj=-0.51 0.16 0.00 instrument_gain_corr=0.00 0.00 0.00 0.00 0.00 0.00" ;
		:Scatterometer\ Processing\ Control = "-limits /sdps/sdpsoper/Science/OCSSW/V2015.2/data/aquarius/scatterometer/L1B_limits_flA_05-08-2012.txt -debug -1 -L2_filter_rfi -param_file /sdps/sdpsoper/Science/OCSSW/V2015.2/data/aquarius/scatterometer/params_pointing_fix_10-31-2012.txt -dir_dat /sdps/sdpsoper/Science/OCSSW/V2015.2/data/aquarius/scatterometer -dir_out /data7/sdpsoper/vdc/vpu6/workbuf -dir_scratch /dev/shm/tmp_76630544 -apc_file /sdps/sdpsoper/Science/OCSSW/V2015.2/data/aquarius/scatterometer/L2_APC_matrix_theory_10-04-2011.txt -cal_level 3 -suppress_tlm_warnings -i /data7/sdpsoper/vdc/vpu6/workbuf/Q2014050173000.L1A_SCI " ;
		:_lastModified = "2015155172225000" ;
		:Conventions = "CF-1.6" ;
		:institution = "NASA/GSFC OBPG" ;
		:Number\ of\ Beams = 3 ;
		:Radiometer\ Polarizations = 4 ;
		:Radiometer\ Subcycles = 12 ;
		:Radiometer\ Signals\ per\ Subcycle = 5 ;
		:Scatterometer\ Polarizations = 6 ;
		:Scatterometer\ Subcycles = 8 ;
		:Start\ Time = "2014050173000992" ;
		:Start\ Year = 2014 ;
		:Start\ Day = 50 ;
		:Start\ Millisec = 63000992 ;
		:End\ Year = 2014 ;
		:End\ Day = 50 ;
		:End\ Millisec = 68879074 ;
		:Node\ Crossing\ Time = "2014050175430000" ;
		:Orbit\ Node\ Longitude = 2.48651f ;
		:Latitude\ Units = "degrees North" ;
		:Longitude\ Units = "degrees East" ;
		:Orbit\ Number = 14496 ;
		:Cycle\ Number = 130 ;
		:Pass\ Number = 100 ;
		:Number\ of\ Blocks = 4083 ;
		:End\ Time = "2014050190759074" ;
		:Percent\ Water = 0.7162888f ;
		:Percent\ RFI = 7.042414f ;
		:Mean\ Solar\ 1415\ MHz\ Flux = 113.75f ;
		:RAD_ANCILLARY_FILE1 = "y2014021912.h5:N2014050_SST_OIV2AV_24h.nc,N2014051_SST_OIV2AV_24h.nc,N201405012_QATM_NCEP_6h.h5,N201405012_QMET_NCEP_6h,N201405012_SWH_NCEP_6h.h5,N201405000_SEAICE_NCEP_24h.hdf,N201405100_SEAICE_NCEP_24h.hdf,N201405000_SALINITY_HYCOM_24h.h5" ;
		:RAD_ANCILLARY_FILE2 = "y2014021918.h5:N2014050_SST_OIV2AV_24h.nc,N2014051_SST_OIV2AV_24h.nc,N201405018_QATM_NCEP_6h.h5,N201405018_QMET_NCEP_6h,N201405018_SWH_NCEP_6h.h5,N201405000_SEAICE_NCEP_24h.hdf,N201405100_SEAICE_NCEP_24h.hdf,N201405000_SALINITY_HYCOM_24h.h5" ;
		:RAD_ANCILLARY_FILE3 = "y2014022000.h5:N2014050_SST_OIV2AV_24h.nc,N2014051_SST_OIV2AV_24h.nc,N201405100_QATM_NCEP_6h.h5,N201405100_QMET_NCEP_6h,N201405100_SWH_NCEP_6h.h5,N201405000_SEAICE_NCEP_24h.hdf,N201405100_SEAICE_NCEP_24h.hdf,N201405000_SALINITY_HYCOM_24h.h5" ;
		:Scatterometer\ Ancillary\ Files = "SEAICEFILE1=N201405000_SEAICE_NCEP_24h.hdf,TECFILE1=N201405000_TEC_IGS_24h.h5,QMETFILE1=N201405012_QMET_NCEP_6h,QMETFILE2=N201405018_QMET_NCEP_6h,QMETFILE3=N201405100_QMET_NCEP_6h" ;
		:Radiometer\ Calibration\ Files = "coeff_loss_V4.txt,coeff_nl.txt" ;
		:Radiometer\ Data\ Tables = "land_tables_V3.6.h5,gain_ice_V3.6.h5,tausq.h5,ocean_reflectance.h5,sun_tables_V3.6.h5,sun_bak_tables.h5,galaxy_wind_tables_V2.0.h5,apc_matrix_may2013_1.h5,land_corr_tables_V3.6.h5,error_tab.h5,deW_harm_coeffs_V9A_MI.h5,sigma0_harm_coeffs_V9A_MI.h5,dtbw_residual_win_sigma_bin_flag_V9_HHH_A.h5,dtbw_residual_win_wav_bin_V9_HHH_A.h5,AQ_SSS_clim_map_testbedV41_2year.h5,dta_gal_symm.h5" ;
		:Scatterometer\ Coefficient\ Files = "atc_prt_convert_v3.txt,ext_temps_constants_convert_v3.txt,scat_temps_convert_v1.txt,radiometer_constants_convert_v2.txt,cmd_gn.dat" ;
		:Delta\ TND\ V\ coefficient = 0.005956746f, 0.00631605f, 0.006228931f ;
		:Delta\ TND\ H\ coefficient = 0.005496748f, 0.005015455f, 0.006067232f ;
		:Radiometer\ Flag\ Limits = "RFI: 15 7 Land: 0.001 0.01 Ice: 0.001 0.01 Wind: 15 20 Temp: 1 3 FluxD: 0.02 0.05 FluxR: 0.02 0.05 Glint: 0.02 0.05 Moon: 0.02 0.05 Gal: 0.02 0.05 RPY: 1 1 5 Flare: 5e-05 0.0001 Tb cons: 0.4 Cold Water: 5 0 TF-TA: -1 -0.3 -1 0.3 Refl 1st Stokes (moon): 0.25 0.5 Refl 1st Stokes (galaxy): 5.6 3.6 (wind): 3" ;
		:Nominal\ Navigation = "TRUE" ;
		:Radiometer\ Offset\ Correction = -0.0242684f, 0.0416904f, -0.05682934f, -0.128805f, -0.08102583f, -0.008495356f ;

group: Aquarius\ Data {
  dimensions:
  	phony_dim_0 = 4083 ;
  	phony_dim_1 = 3 ;
  variables:
  	float Kpc_HH_ant(phony_dim_0, phony_dim_1) ;
  		Kpc_HH_ant:long_name = "Kpc statistical uncertainty for ANT HH NRCS" ;
  		Kpc_HH_ant:valid_min = 0.f ;
  		Kpc_HH_ant:valid_max = 0.f ;
  		Kpc_HH_ant:_FillValue = -999.f ;
  	float Kpc_HH_toa(phony_dim_0, phony_dim_1) ;
  		Kpc_HH_toa:long_name = "Kpc statistical uncertainty for TOA HH NRCS" ;
  		Kpc_HH_toa:valid_min = 0.f ;
  		Kpc_HH_toa:valid_max = 0.f ;
  		Kpc_HH_toa:_FillValue = -999.f ;
  	float Kpc_HV_ant(phony_dim_0, phony_dim_1) ;
  		Kpc_HV_ant:long_name = "Kpc statistical uncertainty for ANT HV NRCS" ;
  		Kpc_HV_ant:valid_min = 0.f ;
  		Kpc_HV_ant:valid_max = 0.f ;
  		Kpc_HV_ant:_FillValue = -999.f ;
  	float Kpc_HV_toa(phony_dim_0, phony_dim_1) ;
  		Kpc_HV_toa:long_name = "Kpc statistical uncertainty for TOA HV NRCS" ;
  		Kpc_HV_toa:valid_min = 0.f ;
  		Kpc_HV_toa:valid_max = 0.f ;
  		Kpc_HV_toa:_FillValue = -999.f ;
  	float Kpc_VH_ant(phony_dim_0, phony_dim_1) ;
  		Kpc_VH_ant:long_name = "Kpc statistical uncertainty for ANT VH NRCS" ;
  		Kpc_VH_ant:valid_min = 0.f ;
  		Kpc_VH_ant:valid_max = 0.f ;
  		Kpc_VH_ant:_FillValue = -999.f ;
  	float Kpc_VH_toa(phony_dim_0, phony_dim_1) ;
  		Kpc_VH_toa:long_name = "Kpc statistical uncertainty for TOA VH NRCS" ;
  		Kpc_VH_toa:valid_min = 0.f ;
  		Kpc_VH_toa:valid_max = 0.f ;
  		Kpc_VH_toa:_FillValue = -999.f ;
  	float Kpc_VV_ant(phony_dim_0, phony_dim_1) ;
  		Kpc_VV_ant:long_name = "Kpc statistical uncertainty for ANT VV NRCS" ;
  		Kpc_VV_ant:valid_min = 0.f ;
  		Kpc_VV_ant:valid_max = 0.f ;
  		Kpc_VV_ant:_FillValue = -999.f ;
  	float Kpc_VV_toa(phony_dim_0, phony_dim_1) ;
  		Kpc_VV_toa:long_name = "Kpc statistical uncertainty for TOA VV NRCS" ;
  		Kpc_VV_toa:valid_min = 0.f ;
  		Kpc_VV_toa:valid_max = 0.f ;
  		Kpc_VV_toa:_FillValue = -999.f ;
  	float Kpc_total(phony_dim_0, phony_dim_1) ;
  		Kpc_total:long_name = "Statistical uncertainty for total power NRCS" ;
  		Kpc_total:valid_min = 0.f ;
  		Kpc_total:valid_max = 0.f ;
  		Kpc_total:_FillValue = -999.f ;
  	float SSS(phony_dim_0, phony_dim_1) ;
  		SSS:long_name = "Sea Surface Salinity" ;
  		SSS:valid_min = 0.f ;
  		SSS:valid_max = 0.f ;
  		SSS:units = "PSU" ;
  		SSS:_FillValue = -9999.f ;
  		SSS:standard_name = "sea_surface_salinity" ;
  	float SSS_nolc(phony_dim_0, phony_dim_1) ;
  		SSS_nolc:long_name = "Sea Surface Salinity (nolc)" ;
  		SSS_nolc:valid_min = 0.f ;
  		SSS_nolc:valid_max = 0.f ;
  		SSS_nolc:units = "PSU" ;
  		SSS_nolc:_FillValue = -9999.f ;
  		SSS_nolc:standard_name = "sea_surface_salinity" ;
  	float SSS_unc_ran(phony_dim_0, phony_dim_1) ;
  		SSS_unc_ran:long_name = "Sea Surface Salinity uncertainty (random)" ;
  		SSS_unc_ran:valid_min = 0.f ;
  		SSS_unc_ran:valid_max = 0.f ;
  		SSS_unc_ran:units = "PSU" ;
  		SSS_unc_ran:_FillValue = -9999.f ;
  	float SSS_unc_sys(phony_dim_0, phony_dim_1) ;
  		SSS_unc_sys:long_name = "Sea Surface Salinity uncertainty (systematic)" ;
  		SSS_unc_sys:valid_min = 0.f ;
  		SSS_unc_sys:valid_max = 0.f ;
  		SSS_unc_sys:units = "PSU" ;
  		SSS_unc_sys:_FillValue = -9999.f ;
  	float anc_SSS(phony_dim_0, phony_dim_1) ;
  		anc_SSS:long_name = "Sea surface salinity (HYCOM)" ;
  		anc_SSS:valid_min = 0.f ;
  		anc_SSS:valid_max = 0.f ;
  		anc_SSS:units = "PSU" ;
  		anc_SSS:_FillValue = -999.f ;
  	float anc_Tb_dw(phony_dim_0, phony_dim_1) ;
  		anc_Tb_dw:long_name = "Downwelling atmospheric brightness temperature" ;
  		anc_Tb_dw:valid_min = 0.f ;
  		anc_Tb_dw:valid_max = 0.f ;
  		anc_Tb_dw:units = "Kelvin" ;
  		anc_Tb_dw:_FillValue = -999.f ;
  	float anc_Tb_up(phony_dim_0, phony_dim_1) ;
  		anc_Tb_up:long_name = "Upwelling atmospheric brightness temperature" ;
  		anc_Tb_up:valid_min = 0.f ;
  		anc_Tb_up:valid_max = 0.f ;
  		anc_Tb_up:units = "Kelvin" ;
  		anc_Tb_up:_FillValue = -999.f ;
  	float anc_cwat(phony_dim_0, phony_dim_1) ;
  		anc_cwat:long_name = "Cloud Water" ;
  		anc_cwat:valid_min = 0.f ;
  		anc_cwat:valid_max = 0.f ;
  		anc_cwat:units = "kg m-2" ;
  		anc_cwat:_FillValue = -999.f ;
  	float anc_sm(phony_dim_0, phony_dim_1) ;
  		anc_sm:long_name = "Soil Moisture" ;
  		anc_sm:valid_min = 0.f ;
  		anc_sm:valid_max = 1.f ;
  		anc_sm:units = "fraction" ;
  		anc_sm:_FillValue = -999.f ;
  	float anc_subsurf_temp(phony_dim_0, phony_dim_1) ;
  		anc_subsurf_temp:long_name = "Sub-Surface Temperature" ;
  		anc_subsurf_temp:valid_min = 0.f ;
  		anc_subsurf_temp:valid_max = 0.f ;
  		anc_subsurf_temp:units = "Kelvin" ;
  		anc_subsurf_temp:_FillValue = -999.f ;
  	float anc_surface_pressure(phony_dim_0, phony_dim_1) ;
  		anc_surface_pressure:long_name = "Surface Pressure" ;
  		anc_surface_pressure:valid_min = 0.f ;
  		anc_surface_pressure:valid_max = 0.f ;
  		anc_surface_pressure:units = "Pascals" ;
  		anc_surface_pressure:_FillValue = -999.f ;
  	float anc_surface_temp(phony_dim_0, phony_dim_1) ;
  		anc_surface_temp:long_name = "Surface Temperature" ;
  		anc_surface_temp:valid_min = 0.f ;
  		anc_surface_temp:valid_max = 0.f ;
  		anc_surface_temp:units = "Kelvin" ;
  		anc_surface_temp:_FillValue = -999.f ;
  	float anc_swe(phony_dim_0, phony_dim_1) ;
  		anc_swe:long_name = "Snow Water Equivalent" ;
  		anc_swe:valid_min = 0.f ;
  		anc_swe:valid_max = 0.f ;
  		anc_swe:units = "kg/m^2" ;
  		anc_swe:_FillValue = -999.f ;
  	float anc_swh(phony_dim_0, phony_dim_1) ;
  		anc_swh:long_name = "Significant wave height" ;
  		anc_swh:valid_min = 0.f ;
  		anc_swh:valid_max = 0.f ;
  		anc_swh:units = "meters" ;
  		anc_swh:_FillValue = -999.f ;
  	float anc_trans(phony_dim_0, phony_dim_1) ;
  		anc_trans:long_name = "Atmospheric Transmittance" ;
  		anc_trans:valid_min = 0.f ;
  		anc_trans:valid_max = 0.f ;
  		anc_trans:_FillValue = -999.f ;
  	float anc_wind_dir(phony_dim_0, phony_dim_1) ;
  		anc_wind_dir:long_name = "Ancillary Wind Direction 10m above surface" ;
  		anc_wind_dir:valid_min = 0.f ;
  		anc_wind_dir:valid_max = 0.f ;
  		anc_wind_dir:units = "degrees" ;
  		anc_wind_dir:_FillValue = -999.f ;
  	float anc_wind_speed(phony_dim_0, phony_dim_1) ;
  		anc_wind_speed:long_name = "Ancillary Wind Speed 10m above surface" ;
  		anc_wind_speed:valid_min = 0.f ;
  		anc_wind_speed:valid_max = 0.f ;
  		anc_wind_speed:units = "meters/sec" ;
  		anc_wind_speed:_FillValue = -999.f ;
  	float density(phony_dim_0, phony_dim_1) ;
  		density:long_name = "Derived Surface Density based on TEOS-10" ;
  		density:valid_min = 0.f ;
  		density:valid_max = 0.f ;
  		density:units = "kg/m^3" ;
  		density:_FillValue = -9999.f ;
  		density:standard_name = "sea_surface_density" ;
  	float rad_Ta3(phony_dim_0, phony_dim_1) ;
  		rad_Ta3:long_name = "Radiometer Ta 3rd Stokes" ;
  		rad_Ta3:valid_min = 0.f ;
  		rad_Ta3:valid_max = 0.f ;
  		rad_Ta3:units = "Kelvin" ;
  		rad_Ta3:_FillValue = -9999.f ;
  	float rad_Ta30(phony_dim_0, phony_dim_1) ;
  		rad_Ta30:long_name = "Radiometer Ta 3rd Stokes (no exp drift)" ;
  		rad_Ta30:valid_max = 0.f ;
  		rad_Ta30:units = "Kelvin" ;
  		rad_Ta30:_FillValue = -9999.f ;
  		rad_Ta30:valid_min = 0.f ;
  	float rad_TaH(phony_dim_0, phony_dim_1) ;
  		rad_TaH:long_name = "Radiometer Ta H polarization" ;
  		rad_TaH:valid_min = 0.f ;
  		rad_TaH:valid_max = 0.f ;
  		rad_TaH:units = "Kelvin" ;
  		rad_TaH:_FillValue = -9999.f ;
  	float rad_TaH0(phony_dim_0, phony_dim_1) ;
  		rad_TaH0:long_name = "Radiometer Ta H polar (no exp drift)" ;
  		rad_TaH0:valid_min = 0.f ;
  		rad_TaH0:valid_max = 0.f ;
  		rad_TaH0:units = "Kelvin" ;
  		rad_TaH0:_FillValue = -9999.f ;
  	float rad_TaV(phony_dim_0, phony_dim_1) ;
  		rad_TaV:long_name = "Radiometer Ta V polarization" ;
  		rad_TaV:valid_min = 0.f ;
  		rad_TaV:valid_max = 0.f ;
  		rad_TaV:units = "Kelvin" ;
  		rad_TaV:_FillValue = -9999.f ;
  	float rad_TaV0(phony_dim_0, phony_dim_1) ;
  		rad_TaV0:long_name = "Radiometer Ta V polar (no exp drift)" ;
  		rad_TaV0:valid_min = 0.f ;
  		rad_TaV0:valid_max = 0.f ;
  		rad_TaV0:units = "Kelvin" ;
  		rad_TaV0:_FillValue = -9999.f ;
  	float rad_TbH(phony_dim_0, phony_dim_1) ;
  		rad_TbH:long_name = "Tb H polarization (no rough corr)" ;
  		rad_TbH:valid_min = 0.f ;
  		rad_TbH:valid_max = 0.f ;
  		rad_TbH:units = "Kelvin" ;
  		rad_TbH:_FillValue = -9999.f ;
  	float rad_TbH_nolc(phony_dim_0, phony_dim_1) ;
  		rad_TbH_nolc:long_name = "Earth surface Tb H polarization (nolc)" ;
  		rad_TbH_nolc:valid_min = 0.f ;
  		rad_TbH_nolc:valid_max = 0.f ;
  		rad_TbH_nolc:units = "Kelvin" ;
  		rad_TbH_nolc:_FillValue = -9999.f ;
  	float rad_TbH_rc(phony_dim_0, phony_dim_1) ;
  		rad_TbH_rc:long_name = "Tb H polarization (rough corr)" ;
  		rad_TbH_rc:valid_min = 0.f ;
  		rad_TbH_rc:valid_max = 0.f ;
  		rad_TbH_rc:units = "Kelvin" ;
  		rad_TbH_rc:_FillValue = -9999.f ;
  	float rad_TbH_rc_nolc(phony_dim_0, phony_dim_1) ;
  		rad_TbH_rc_nolc:long_name = "Tb H polarization (roughness corr, nolc)" ;
  		rad_TbH_rc_nolc:valid_min = 0.f ;
  		rad_TbH_rc_nolc:valid_max = 0.f ;
  		rad_TbH_rc_nolc:units = "Kelvin" ;
  		rad_TbH_rc_nolc:_FillValue = -9999.f ;
  	float rad_TbV(phony_dim_0, phony_dim_1) ;
  		rad_TbV:long_name = "Tb V polarization (no rough corr)" ;
  		rad_TbV:valid_min = 0.f ;
  		rad_TbV:valid_max = 0.f ;
  		rad_TbV:units = "Kelvin" ;
  		rad_TbV:_FillValue = -9999.f ;
  	float rad_TbV_nolc(phony_dim_0, phony_dim_1) ;
  		rad_TbV_nolc:long_name = "Earth surface Tb V polarization (no lc)" ;
  		rad_TbV_nolc:valid_min = 0.f ;
  		rad_TbV_nolc:valid_max = 0.f ;
  		rad_TbV_nolc:units = "Kelvin" ;
  		rad_TbV_nolc:_FillValue = -9999.f ;
  	float rad_TbV_rc(phony_dim_0, phony_dim_1) ;
  		rad_TbV_rc:long_name = "Tb V polarization (rough corr)" ;
  		rad_TbV_rc:valid_min = 0.f ;
  		rad_TbV_rc:valid_max = 0.f ;
  		rad_TbV_rc:units = "Kelvin" ;
  		rad_TbV_rc:_FillValue = -9999.f ;
  	float rad_TbV_rc_nolc(phony_dim_0, phony_dim_1) ;
  		rad_TbV_rc_nolc:long_name = "Tb V polarization (roughness corr, nolc)" ;
  		rad_TbV_rc_nolc:valid_min = 0.f ;
  		rad_TbV_rc_nolc:valid_max = 0.f ;
  		rad_TbV_rc_nolc:units = "Kelvin" ;
  		rad_TbV_rc_nolc:_FillValue = -9999.f ;
  	float rad_Tb_consistency(phony_dim_0, phony_dim_1) ;
  		rad_Tb_consistency:long_name = "Tb consistency check" ;
  		rad_Tb_consistency:valid_min = 0.f ;
  		rad_Tb_consistency:valid_max = 0.f ;
  		rad_Tb_consistency:units = "Kelvin" ;
  		rad_Tb_consistency:_FillValue = -9999.f ;
  	float rad_Tb_consistency_nolc(phony_dim_0, phony_dim_1) ;
  		rad_Tb_consistency_nolc:long_name = "Tb consistency check (nolc)" ;
  		rad_Tb_consistency_nolc:valid_min = 0.f ;
  		rad_Tb_consistency_nolc:valid_max = 0.f ;
  		rad_Tb_consistency_nolc:units = "Kelvin" ;
  		rad_Tb_consistency_nolc:_FillValue = -9999.f ;
  	float rad_Tf3(phony_dim_0, phony_dim_1) ;
  		rad_Tf3:long_name = "Radiometer Ta 3rd Stokes (rfi filtered)" ;
  		rad_Tf3:valid_min = 0.f ;
  		rad_Tf3:valid_max = 0.f ;
  		rad_Tf3:units = "Kelvin" ;
  		rad_Tf3:_FillValue = -9999.f ;
  	float rad_Tf30(phony_dim_0, phony_dim_1) ;
  		rad_Tf30:long_name = "Radiometer Ta 3 (rfi filtered/no exp drift)" ;
  		rad_Tf30:valid_min = 0.f ;
  		rad_Tf30:valid_max = 0.f ;
  		rad_Tf30:units = "Kelvin" ;
  		rad_Tf30:_FillValue = -9999.f ;
  	float rad_TfH(phony_dim_0, phony_dim_1) ;
  		rad_TfH:long_name = "Radiometer Ta H polarization (rfi filtered)" ;
  		rad_TfH:valid_min = 0.f ;
  		rad_TfH:valid_max = 0.f ;
  		rad_TfH:units = "Kelvin" ;
  		rad_TfH:_FillValue = -9999.f ;
  	float rad_TfH0(phony_dim_0, phony_dim_1) ;
  		rad_TfH0:long_name = "Radiometer Ta H (rfi filtered/no exp drift)" ;
  		rad_TfH0:valid_min = 0.f ;
  		rad_TfH0:valid_max = 0.f ;
  		rad_TfH0:units = "Kelvin" ;
  		rad_TfH0:_FillValue = -9999.f ;
  	float rad_TfV(phony_dim_0, phony_dim_1) ;
  		rad_TfV:long_name = "Radiometer Ta V polarization (rfi filtered)" ;
  		rad_TfV:valid_min = 0.f ;
  		rad_TfV:valid_max = 0.f ;
  		rad_TfV:units = "Kelvin" ;
  		rad_TfV:_FillValue = -9999.f ;
  	float rad_TfV0(phony_dim_0, phony_dim_1) ;
  		rad_TfV0:long_name = "Radiometer Ta V (rfi filtered/no exp drift)" ;
  		rad_TfV0:valid_min = 0.f ;
  		rad_TfV0:valid_max = 0.f ;
  		rad_TfV0:units = "Kelvin" ;
  		rad_TfV0:_FillValue = -9999.f ;
  	float rad_dtb_sst_wspd_H(phony_dim_0, phony_dim_1) ;
  		rad_dtb_sst_wspd_H:long_name = "Radiometer SST bias emissivity correction H" ;
  		rad_dtb_sst_wspd_H:valid_min = 0.f ;
  		rad_dtb_sst_wspd_H:valid_max = 0.f ;
  		rad_dtb_sst_wspd_H:units = "Kelvin" ;
  		rad_dtb_sst_wspd_H:_FillValue = -9999.f ;
  	float rad_dtb_sst_wspd_V(phony_dim_0, phony_dim_1) ;
  		rad_dtb_sst_wspd_V:long_name = "Radiometer SST bias emissivity correction V" ;
  		rad_dtb_sst_wspd_V:valid_min = 0.f ;
  		rad_dtb_sst_wspd_V:valid_max = 0.f ;
  		rad_dtb_sst_wspd_V:units = "Kelvin" ;
  		rad_dtb_sst_wspd_V:_FillValue = -9999.f ;
  	float rad_exp_Ta3(phony_dim_0, phony_dim_1) ;
  		rad_exp_Ta3:long_name = "Radiometer Ta 3rd Stokes (expected)" ;
  		rad_exp_Ta3:valid_min = 0.f ;
  		rad_exp_Ta3:valid_max = 0.f ;
  		rad_exp_Ta3:units = "Kelvin" ;
  		rad_exp_Ta3:_FillValue = -9999.f ;
  	float rad_exp_Ta3_hhh(phony_dim_0, phony_dim_1) ;
  		rad_exp_Ta3_hhh:long_name = "Radiometer Ta 3rd Stokes (expected/HHH winds)" ;
  		rad_exp_Ta3_hhh:valid_min = 0.f ;
  		rad_exp_Ta3_hhh:valid_max = 0.f ;
  		rad_exp_Ta3_hhh:units = "Kelvin" ;
  		rad_exp_Ta3_hhh:_FillValue = -9999.f ;
  	float rad_exp_TaH(phony_dim_0, phony_dim_1) ;
  		rad_exp_TaH:long_name = "Radiometer Ta H (expected)" ;
  		rad_exp_TaH:valid_min = 0.f ;
  		rad_exp_TaH:valid_max = 0.f ;
  		rad_exp_TaH:units = "Kelvin" ;
  		rad_exp_TaH:_FillValue = -9999.f ;
  	float rad_exp_TaH_hhh(phony_dim_0, phony_dim_1) ;
  		rad_exp_TaH_hhh:long_name = "Radiometer Ta H (expected/HHH winds)" ;
  		rad_exp_TaH_hhh:valid_min = 0.f ;
  		rad_exp_TaH_hhh:valid_max = 0.f ;
  		rad_exp_TaH_hhh:units = "Kelvin" ;
  		rad_exp_TaH_hhh:_FillValue = -9999.f ;
  	float rad_exp_TaV(phony_dim_0, phony_dim_1) ;
  		rad_exp_TaV:long_name = "Radiometer Ta V (expected)" ;
  		rad_exp_TaV:valid_min = 0.f ;
  		rad_exp_TaV:valid_max = 0.f ;
  		rad_exp_TaV:units = "Kelvin" ;
  		rad_exp_TaV:_FillValue = -9999.f ;
  	float rad_exp_TaV_hhh(phony_dim_0, phony_dim_1) ;
  		rad_exp_TaV_hhh:long_name = "Radiometer Ta V (expected/HHH winds)" ;
  		rad_exp_TaV_hhh:valid_min = 0.f ;
  		rad_exp_TaV_hhh:valid_max = 0.f ;
  		rad_exp_TaV_hhh:units = "Kelvin" ;
  		rad_exp_TaV_hhh:_FillValue = -9999.f ;
  	float rad_exp_TbH(phony_dim_0, phony_dim_1) ;
  		rad_exp_TbH:long_name = "Radiometer Tb H (expected)" ;
  		rad_exp_TbH:valid_min = 0.f ;
  		rad_exp_TbH:valid_max = 0.f ;
  		rad_exp_TbH:units = "Kelvin" ;
  		rad_exp_TbH:_FillValue = -9999.f ;
  	float rad_exp_TbH0(phony_dim_0, phony_dim_1) ;
  		rad_exp_TbH0:long_name = "Radiometer Tb H (expected smooth)" ;
  		rad_exp_TbH0:valid_min = 0.f ;
  		rad_exp_TbH0:valid_max = 0.f ;
  		rad_exp_TbH0:units = "Kelvin" ;
  		rad_exp_TbH0:_FillValue = -9999.f ;
  	float rad_exp_TbV(phony_dim_0, phony_dim_1) ;
  		rad_exp_TbV:long_name = "Radiometer Tb V (expected)" ;
  		rad_exp_TbV:valid_min = 0.f ;
  		rad_exp_TbV:valid_max = 0.f ;
  		rad_exp_TbV:units = "Kelvin" ;
  		rad_exp_TbV:_FillValue = -9999.f ;
  	float rad_exp_TbV0(phony_dim_0, phony_dim_1) ;
  		rad_exp_TbV0:long_name = "Radiometer Tb V (expected smooth)" ;
  		rad_exp_TbV0:valid_min = 0.f ;
  		rad_exp_TbV0:valid_max = 0.f ;
  		rad_exp_TbV0:units = "Kelvin" ;
  		rad_exp_TbV0:_FillValue = -9999.f ;
  	float rad_far_TaH(phony_dim_0, phony_dim_1) ;
  		rad_far_TaH:long_name = "Radiometer Faraday Angle" ;
  		rad_far_TaH:valid_min = 0.f ;
  		rad_far_TaH:valid_max = 0.f ;
  		rad_far_TaH:units = "Degrees" ;
  		rad_far_TaH:_FillValue = -9999.f ;
  	float rad_galact_Ta_dir_3(phony_dim_0, phony_dim_1) ;
  		rad_galact_Ta_dir_3:long_name = "Radiometer Galactic Direct Corr 3rd Stokes" ;
  		rad_galact_Ta_dir_3:valid_min = 0.f ;
  		rad_galact_Ta_dir_3:valid_max = 0.f ;
  		rad_galact_Ta_dir_3:units = "Kelvin" ;
  		rad_galact_Ta_dir_3:_FillValue = -9999.f ;
  	float rad_galact_Ta_dir_H(phony_dim_0, phony_dim_1) ;
  		rad_galact_Ta_dir_H:long_name = "Radiometer Galactic Direct Corr H polar" ;
  		rad_galact_Ta_dir_H:valid_min = 0.f ;
  		rad_galact_Ta_dir_H:valid_max = 0.f ;
  		rad_galact_Ta_dir_H:units = "Kelvin" ;
  		rad_galact_Ta_dir_H:_FillValue = -9999.f ;
  	float rad_galact_Ta_dir_V(phony_dim_0, phony_dim_1) ;
  		rad_galact_Ta_dir_V:long_name = "Radiometer Galactic Direct Corr V polar" ;
  		rad_galact_Ta_dir_V:valid_min = 0.f ;
  		rad_galact_Ta_dir_V:valid_max = 0.f ;
  		rad_galact_Ta_dir_V:units = "Kelvin" ;
  		rad_galact_Ta_dir_V:_FillValue = -9999.f ;
  	float rad_galact_Ta_ref_3(phony_dim_0, phony_dim_1) ;
  		rad_galact_Ta_ref_3:long_name = "Radiometer Galactic Reflect Corr 3rd Stokes" ;
  		rad_galact_Ta_ref_3:valid_min = 0.f ;
  		rad_galact_Ta_ref_3:valid_max = 0.f ;
  		rad_galact_Ta_ref_3:units = "Kelvin" ;
  		rad_galact_Ta_ref_3:_FillValue = -9999.f ;
  	float rad_galact_Ta_ref_GO_H(phony_dim_0, phony_dim_1) ;
  		rad_galact_Ta_ref_GO_H:long_name = "Radiometer Gal Reflect Corr H polar (GO)" ;
  		rad_galact_Ta_ref_GO_H:valid_min = 0.f ;
  		rad_galact_Ta_ref_GO_H:valid_max = 0.f ;
  		rad_galact_Ta_ref_GO_H:units = "Kelvin" ;
  		rad_galact_Ta_ref_GO_H:_FillValue = -9999.f ;
  	float rad_galact_Ta_ref_GO_V(phony_dim_0, phony_dim_1) ;
  		rad_galact_Ta_ref_GO_V:long_name = "Radiometer Gal Reflect Corr V polar (GO)" ;
  		rad_galact_Ta_ref_GO_V:valid_min = 0.f ;
  		rad_galact_Ta_ref_GO_V:valid_max = 0.f ;
  		rad_galact_Ta_ref_GO_V:units = "Kelvin" ;
  		rad_galact_Ta_ref_GO_V:_FillValue = -9999.f ;
  	float rad_galact_Ta_ref_H(phony_dim_0, phony_dim_1) ;
  		rad_galact_Ta_ref_H:long_name = "Radiometer Galactic Reflect Corr H polar" ;
  		rad_galact_Ta_ref_H:valid_min = 0.f ;
  		rad_galact_Ta_ref_H:valid_max = 0.f ;
  		rad_galact_Ta_ref_H:units = "Kelvin" ;
  		rad_galact_Ta_ref_H:_FillValue = -9999.f ;
  	float rad_galact_Ta_ref_V(phony_dim_0, phony_dim_1) ;
  		rad_galact_Ta_ref_V:long_name = "Radiometer Galactic Reflect Corr V polar" ;
  		rad_galact_Ta_ref_V:valid_min = 0.f ;
  		rad_galact_Ta_ref_V:valid_max = 0.f ;
  		rad_galact_Ta_ref_V:units = "Kelvin" ;
  		rad_galact_Ta_ref_V:_FillValue = -9999.f ;
  	float rad_galact_dTa_H(phony_dim_0, phony_dim_1) ;
  		rad_galact_dTa_H:long_name = "Empirical Gal Reflect Adj H polar" ;
  		rad_galact_dTa_H:valid_min = 0.f ;
  		rad_galact_dTa_H:valid_max = 0.f ;
  		rad_galact_dTa_H:units = "Kelvin" ;
  		rad_galact_dTa_H:_FillValue = -9999.f ;
  	float rad_galact_dTa_V(phony_dim_0, phony_dim_1) ;
  		rad_galact_dTa_V:long_name = "Empirical Gal Reflect Adj V polar" ;
  		rad_galact_dTa_V:valid_min = 0.f ;
  		rad_galact_dTa_V:valid_max = 0.f ;
  		rad_galact_dTa_V:units = "Kelvin" ;
  		rad_galact_dTa_V:_FillValue = -9999.f ;
  	float rad_hh_wind_speed(phony_dim_0, phony_dim_1) ;
  		rad_hh_wind_speed:long_name = "Radiometer HH wind speed" ;
  		rad_hh_wind_speed:valid_min = 0.f ;
  		rad_hh_wind_speed:valid_max = 0.f ;
  		rad_hh_wind_speed:units = "meters/sec" ;
  		rad_hh_wind_speed:_FillValue = -9999.f ;
  	float rad_hhh_wind_speed(phony_dim_0, phony_dim_1) ;
  		rad_hhh_wind_speed:long_name = "Radiometer HHH wind speed" ;
  		rad_hhh_wind_speed:valid_min = 0.f ;
  		rad_hhh_wind_speed:valid_max = 0.f ;
  		rad_hhh_wind_speed:units = "meters/sec" ;
  		rad_hhh_wind_speed:_FillValue = -9999.f ;
  	float rad_ice_frac(phony_dim_0, phony_dim_1) ;
  		rad_ice_frac:long_name = "Fraction of ice contamination (radiometer)" ;
  		rad_ice_frac:valid_min = 0.f ;
  		rad_ice_frac:valid_max = 0.f ;
  		rad_ice_frac:_FillValue = -9999.f ;
  	float rad_land_frac(phony_dim_0, phony_dim_1) ;
  		rad_land_frac:long_name = "Fraction of land contamination (radiometer)" ;
  		rad_land_frac:valid_min = 0.f ;
  		rad_land_frac:valid_max = 0.f ;
  		rad_land_frac:_FillValue = -9999.f ;
  	float rad_moon_Ta_ref_3(phony_dim_0, phony_dim_1) ;
  		rad_moon_Ta_ref_3:long_name = "Radiometer Lunar Reflect Corr 3rd Stokes" ;
  		rad_moon_Ta_ref_3:valid_min = 0.f ;
  		rad_moon_Ta_ref_3:valid_max = 0.f ;
  		rad_moon_Ta_ref_3:units = "Kelvin" ;
  		rad_moon_Ta_ref_3:_FillValue = -9999.f ;
  	float rad_moon_Ta_ref_H(phony_dim_0, phony_dim_1) ;
  		rad_moon_Ta_ref_H:long_name = "Radiometer Lunar Reflect Corr H polar" ;
  		rad_moon_Ta_ref_H:valid_min = 0.f ;
  		rad_moon_Ta_ref_H:valid_max = 0.f ;
  		rad_moon_Ta_ref_H:units = "Kelvin" ;
  		rad_moon_Ta_ref_H:_FillValue = -9999.f ;
  	float rad_moon_Ta_ref_V(phony_dim_0, phony_dim_1) ;
  		rad_moon_Ta_ref_V:long_name = "Radiometer Lunar Reflect Corr V polar" ;
  		rad_moon_Ta_ref_V:valid_min = 0.f ;
  		rad_moon_Ta_ref_V:valid_max = 0.f ;
  		rad_moon_Ta_ref_V:units = "Kelvin" ;
  		rad_moon_Ta_ref_V:_FillValue = -9999.f ;
  	float rad_solar_Ta_bak_3(phony_dim_0, phony_dim_1) ;
  		rad_solar_Ta_bak_3:long_name = "Radiometer Solar Back Scattered 3rd Stokes" ;
  		rad_solar_Ta_bak_3:valid_min = 0.f ;
  		rad_solar_Ta_bak_3:valid_max = 0.f ;
  		rad_solar_Ta_bak_3:units = "Kelvin" ;
  		rad_solar_Ta_bak_3:_FillValue = -9999.f ;
  	float rad_solar_Ta_bak_H(phony_dim_0, phony_dim_1) ;
  		rad_solar_Ta_bak_H:long_name = "Radiometer Solar Back Scattered H polar" ;
  		rad_solar_Ta_bak_H:valid_min = 0.f ;
  		rad_solar_Ta_bak_H:valid_max = 0.f ;
  		rad_solar_Ta_bak_H:units = "Kelvin" ;
  		rad_solar_Ta_bak_H:_FillValue = -9999.f ;
  	float rad_solar_Ta_bak_V(phony_dim_0, phony_dim_1) ;
  		rad_solar_Ta_bak_V:long_name = "Radiometer Solar Back Scattered V polar" ;
  		rad_solar_Ta_bak_V:valid_min = 0.f ;
  		rad_solar_Ta_bak_V:valid_max = 0.f ;
  		rad_solar_Ta_bak_V:units = "Kelvin" ;
  		rad_solar_Ta_bak_V:_FillValue = -9999.f ;
  	float rad_solar_Ta_dir_3(phony_dim_0, phony_dim_1) ;
  		rad_solar_Ta_dir_3:long_name = "Radiometer Solar Direct Corr 3rd Stokes" ;
  		rad_solar_Ta_dir_3:valid_min = 0.f ;
  		rad_solar_Ta_dir_3:valid_max = 0.f ;
  		rad_solar_Ta_dir_3:units = "Kelvin" ;
  		rad_solar_Ta_dir_3:_FillValue = -9999.f ;
  	float rad_solar_Ta_dir_H(phony_dim_0, phony_dim_1) ;
  		rad_solar_Ta_dir_H:long_name = "Radiometer Solar Direct Corr H polar" ;
  		rad_solar_Ta_dir_H:valid_min = 0.f ;
  		rad_solar_Ta_dir_H:valid_max = 0.f ;
  		rad_solar_Ta_dir_H:units = "Kelvin" ;
  		rad_solar_Ta_dir_H:_FillValue = -9999.f ;
  	float rad_solar_Ta_dir_V(phony_dim_0, phony_dim_1) ;
  		rad_solar_Ta_dir_V:long_name = "Radiometer Solar Direct Corr V polar" ;
  		rad_solar_Ta_dir_V:valid_min = 0.f ;
  		rad_solar_Ta_dir_V:valid_max = 0.f ;
  		rad_solar_Ta_dir_V:units = "Kelvin" ;
  		rad_solar_Ta_dir_V:_FillValue = -9999.f ;
  	float rad_solar_Ta_ref_3(phony_dim_0, phony_dim_1) ;
  		rad_solar_Ta_ref_3:long_name = "Radiometer Solar Reflect Corr 3rd Stokes" ;
  		rad_solar_Ta_ref_3:valid_min = 0.f ;
  		rad_solar_Ta_ref_3:valid_max = 0.f ;
  		rad_solar_Ta_ref_3:units = "Kelvin" ;
  		rad_solar_Ta_ref_3:_FillValue = -9999.f ;
  	float rad_solar_Ta_ref_H(phony_dim_0, phony_dim_1) ;
  		rad_solar_Ta_ref_H:long_name = "Radiometer Solar Reflect Corr H polar" ;
  		rad_solar_Ta_ref_H:valid_min = 0.f ;
  		rad_solar_Ta_ref_H:valid_max = 0.f ;
  		rad_solar_Ta_ref_H:units = "Kelvin" ;
  		rad_solar_Ta_ref_H:_FillValue = -9999.f ;
  	float rad_solar_Ta_ref_V(phony_dim_0, phony_dim_1) ;
  		rad_solar_Ta_ref_V:long_name = "Radiometer Solar Reflect Corr V polar" ;
  		rad_solar_Ta_ref_V:valid_min = 0.f ;
  		rad_solar_Ta_ref_V:valid_max = 0.f ;
  		rad_solar_Ta_ref_V:units = "Kelvin" ;
  		rad_solar_Ta_ref_V:_FillValue = -9999.f ;
  	float rad_toa_H(phony_dim_0, phony_dim_1) ;
  		rad_toa_H:long_name = "Radiometer TOA Tb H polarization" ;
  		rad_toa_H:valid_min = 0.f ;
  		rad_toa_H:valid_max = 0.f ;
  		rad_toa_H:units = "Kelvin" ;
  		rad_toa_H:_FillValue = -9999.f ;
  	float rad_toa_H_nolc(phony_dim_0, phony_dim_1) ;
  		rad_toa_H_nolc:long_name = "Radiometer TOA Tb H polarization (nolc)" ;
  		rad_toa_H_nolc:valid_min = 0.f ;
  		rad_toa_H_nolc:valid_max = 0.f ;
  		rad_toa_H_nolc:units = "Kelvin" ;
  		rad_toa_H_nolc:_FillValue = -9999.f ;
  	float rad_toa_V(phony_dim_0, phony_dim_1) ;
  		rad_toa_V:long_name = "Radiometer TOA Tb V polarization" ;
  		rad_toa_V:valid_min = 0.f ;
  		rad_toa_V:valid_max = 0.f ;
  		rad_toa_V:units = "Kelvin" ;
  		rad_toa_V:_FillValue = -9999.f ;
  	float rad_toa_V_nolc(phony_dim_0, phony_dim_1) ;
  		rad_toa_V_nolc:long_name = "Radiometer TOA Tb V polarization (nolc)" ;
  		rad_toa_V_nolc:valid_min = 0.f ;
  		rad_toa_V_nolc:valid_max = 0.f ;
  		rad_toa_V_nolc:units = "Kelvin" ;
  		rad_toa_V_nolc:_FillValue = -9999.f ;
  	float rad_toi_3(phony_dim_0, phony_dim_1) ;
  		rad_toi_3:long_name = "Radiometer TOI Tb 3rd Stokes" ;
  		rad_toi_3:valid_min = 0.f ;
  		rad_toi_3:valid_max = 0.f ;
  		rad_toi_3:units = "Kelvin" ;
  		rad_toi_3:_FillValue = -9999.f ;
  	float rad_toi_H(phony_dim_0, phony_dim_1) ;
  		rad_toi_H:long_name = "Radiometer TOI Tb H polarization" ;
  		rad_toi_H:valid_min = 0.f ;
  		rad_toi_H:valid_max = 0.f ;
  		rad_toi_H:units = "Kelvin" ;
  		rad_toi_H:_FillValue = -9999.f ;
  	float rad_toi_V(phony_dim_0, phony_dim_1) ;
  		rad_toi_V:long_name = "Radiometer TOI Tb V polarization" ;
  		rad_toi_V:units = "Kelvin" ;
  		rad_toi_V:_FillValue = -9999.f ;
  		rad_toi_V:valid_min = 0.f ;
  		rad_toi_V:valid_max = 0.f ;
  	float scat_HH_ant(phony_dim_0, phony_dim_1) ;
  		scat_HH_ant:long_name = "ANT Scatterometer NRCS for HH polarization" ;
  		scat_HH_ant:valid_min = 0.f ;
  		scat_HH_ant:valid_max = 0.f ;
  		scat_HH_ant:units = "db" ;
  		scat_HH_ant:_FillValue = -999.f ;
  	float scat_HH_exp(phony_dim_0, phony_dim_1) ;
  		scat_HH_exp:long_name = "Expected Sigma0 for HH polarization" ;
  		scat_HH_exp:valid_min = 0.f ;
  		scat_HH_exp:valid_max = 0.f ;
  		scat_HH_exp:units = "db" ;
  		scat_HH_exp:_FillValue = -999.f ;
  	float scat_HH_toa(phony_dim_0, phony_dim_1) ;
  		scat_HH_toa:long_name = "TOA Scatterometer NRCS for HH polarization" ;
  		scat_HH_toa:valid_min = 0.f ;
  		scat_HH_toa:valid_max = 0.f ;
  		scat_HH_toa:units = "db" ;
  		scat_HH_toa:_FillValue = -999.f ;
  	float scat_HV_ant(phony_dim_0, phony_dim_1) ;
  		scat_HV_ant:long_name = "ANT Scatterometer NRCS for HV polarization" ;
  		scat_HV_ant:valid_min = 0.f ;
  		scat_HV_ant:valid_max = 0.f ;
  		scat_HV_ant:units = "db" ;
  		scat_HV_ant:_FillValue = -999.f ;
  	float scat_HV_exp(phony_dim_0, phony_dim_1) ;
  		scat_HV_exp:long_name = "Expected Sigma0 for HV polarization" ;
  		scat_HV_exp:valid_min = 0.f ;
  		scat_HV_exp:valid_max = 0.f ;
  		scat_HV_exp:units = "db" ;
  		scat_HV_exp:_FillValue = -999.f ;
  	float scat_HV_toa(phony_dim_0, phony_dim_1) ;
  		scat_HV_toa:long_name = "TOA Scatterometer NRCS for HV polarization" ;
  		scat_HV_toa:valid_min = 0.f ;
  		scat_HV_toa:valid_max = 0.f ;
  		scat_HV_toa:units = "db" ;
  		scat_HV_toa:_FillValue = -999.f ;
  	float scat_VH_ant(phony_dim_0, phony_dim_1) ;
  		scat_VH_ant:long_name = "ANT Scatterometer NRCS for VH polarization" ;
  		scat_VH_ant:valid_min = 0.f ;
  		scat_VH_ant:valid_max = 0.f ;
  		scat_VH_ant:units = "db" ;
  		scat_VH_ant:_FillValue = -999.f ;
  	float scat_VH_exp(phony_dim_0, phony_dim_1) ;
  		scat_VH_exp:long_name = "Expected Sigma0 for VH polarization" ;
  		scat_VH_exp:valid_min = 0.f ;
  		scat_VH_exp:valid_max = 0.f ;
  		scat_VH_exp:units = "db" ;
  		scat_VH_exp:_FillValue = -999.f ;
  	float scat_VH_toa(phony_dim_0, phony_dim_1) ;
  		scat_VH_toa:long_name = "TOA Scatterometer NRCS for VH polarization" ;
  		scat_VH_toa:valid_min = 0.f ;
  		scat_VH_toa:valid_max = 0.f ;
  		scat_VH_toa:units = "db" ;
  		scat_VH_toa:_FillValue = -999.f ;
  	float scat_VV_ant(phony_dim_0, phony_dim_1) ;
  		scat_VV_ant:long_name = "ANT Scatterometer NRCS for VV polarization" ;
  		scat_VV_ant:valid_min = 0.f ;
  		scat_VV_ant:valid_max = 0.f ;
  		scat_VV_ant:units = "db" ;
  		scat_VV_ant:_FillValue = -999.f ;
  	float scat_VV_exp(phony_dim_0, phony_dim_1) ;
  		scat_VV_exp:long_name = "Expected Sigma0 for VV polarization" ;
  		scat_VV_exp:valid_min = 0.f ;
  		scat_VV_exp:valid_max = 0.f ;
  		scat_VV_exp:units = "db" ;
  		scat_VV_exp:_FillValue = -999.f ;
  	float scat_VV_toa(phony_dim_0, phony_dim_1) ;
  		scat_VV_toa:long_name = "TOA Scatterometer NRCS for VV polarization" ;
  		scat_VV_toa:valid_min = 0.f ;
  		scat_VV_toa:valid_max = 0.f ;
  		scat_VV_toa:units = "db" ;
  		scat_VV_toa:_FillValue = -999.f ;
  	float scat_esurf_H(phony_dim_0, phony_dim_1) ;
  		scat_esurf_H:long_name = "excess surface scatterometer emissivity (H pol)" ;
  		scat_esurf_H:valid_min = 0.f ;
  		scat_esurf_H:valid_max = 0.f ;
  		scat_esurf_H:units = "Kelvin" ;
  		scat_esurf_H:_FillValue = -999.f ;
  	float scat_esurf_H_uncertainty(phony_dim_0, phony_dim_1) ;
  		scat_esurf_H_uncertainty:long_name = "Uncertainty in surface emmissivity (H-pol)" ;
  		scat_esurf_H_uncertainty:valid_min = 0.f ;
  		scat_esurf_H_uncertainty:valid_max = 0.f ;
  		scat_esurf_H_uncertainty:units = "Kelvin" ;
  		scat_esurf_H_uncertainty:_FillValue = -999.f ;
  	float scat_esurf_V(phony_dim_0, phony_dim_1) ;
  		scat_esurf_V:long_name = "excess surface scatterometer emissivity (V pol)" ;
  		scat_esurf_V:valid_min = 0.f ;
  		scat_esurf_V:valid_max = 0.f ;
  		scat_esurf_V:units = "Kelvin" ;
  		scat_esurf_V:_FillValue = -999.f ;
  	float scat_esurf_V_uncertainty(phony_dim_0, phony_dim_1) ;
  		scat_esurf_V_uncertainty:long_name = "Uncertainty in surface emmissivity (V-pol)" ;
  		scat_esurf_V_uncertainty:valid_min = 0.f ;
  		scat_esurf_V_uncertainty:valid_max = 0.f ;
  		scat_esurf_V_uncertainty:units = "Kelvin" ;
  		scat_esurf_V_uncertainty:_FillValue = -999.f ;
  	float scat_ice_frac(phony_dim_0, phony_dim_1) ;
  		scat_ice_frac:long_name = "Fraction of ice contamination (scatterometer)" ;
  		scat_ice_frac:valid_min = 0.f ;
  		scat_ice_frac:valid_max = 0.f ;
  		scat_ice_frac:_FillValue = -999.f ;
  	float scat_land_frac(phony_dim_0, phony_dim_1) ;
  		scat_land_frac:long_name = "Fraction of land contamination (scatterometer)" ;
  		scat_land_frac:valid_min = 0.f ;
  		scat_land_frac:valid_max = 0.f ;
  		scat_land_frac:_FillValue = -999.f ;
  	float scat_tot_toa(phony_dim_0, phony_dim_1) ;
  		scat_tot_toa:long_name = "TOA Scatterometer (Total)" ;
  		scat_tot_toa:valid_min = 0.f ;
  		scat_tot_toa:valid_max = 0.f ;
  		scat_tot_toa:units = "db" ;
  		scat_tot_toa:_FillValue = -999.f ;
  	float scat_wind_speed(phony_dim_0, phony_dim_1) ;
  		scat_wind_speed:long_name = "Scatterometer Wind Speed" ;
  		scat_wind_speed:valid_max = 0.f ;
  		scat_wind_speed:units = "meters/sec" ;
  		scat_wind_speed:_FillValue = -999.f ;
  		scat_wind_speed:valid_min = 0.f ;
  	float wind_uncertainty(phony_dim_0, phony_dim_1) ;
  		wind_uncertainty:long_name = "Estimated wind speed error" ;
  		wind_uncertainty:valid_min = 0.f ;
  		wind_uncertainty:valid_max = 0.f ;
  		wind_uncertainty:units = "meters/sec" ;
  		wind_uncertainty:_FillValue = -999.f ;
  } // group Aquarius\ Data

group: Aquarius\ Flags {
  dimensions:
  	phony_dim_2 = 4083 ;
  	phony_dim_3 = 3 ;
  	phony_dim_4 = 4 ;
  	phony_dim_5 = 12 ;
  	phony_dim_6 = 2 ;
  variables:
  	ubyte rad_rfi_flags(phony_dim_2, phony_dim_3, phony_dim_4, phony_dim_5) ;
  		rad_rfi_flags:long_name = "Radiometer RFI flags" ;
  		rad_rfi_flags:valid_min = 0UB ;
  		rad_rfi_flags:valid_max = 0UB ;
  	uint radiometer_flags(phony_dim_2, phony_dim_3, phony_dim_4) ;
  		radiometer_flags:long_name = "Radiometer data quality flags" ;
  		radiometer_flags:RFI\ contamination = "RFI" ;
  		radiometer_flags:Rain\ in\ main\ beam = "RAIN" ;
  		radiometer_flags:Land\ contamination = "LAND" ;
  		radiometer_flags:Sea\ ice\ contamination = "ICE" ;
  		radiometer_flags:Wind/foam\ contamination = "WIND" ;
  		radiometer_flags:Unusual\ brighness\ temperature = "TEMP" ;
  		radiometer_flags:Direct\ solar\ flux\ contamination = "FLUXD" ;
  		radiometer_flags:Reflected\ solar\ flux\ contamination = "FLUXR" ;
  		radiometer_flags:Sun\ glint = "SUNGLINT" ;
  		radiometer_flags:Moon\ contamination = "MOON" ;
  		radiometer_flags:Galactic\ contamination = "GALACTIC" ;
  		radiometer_flags:Non-nominal\ navigation = "NAV" ;
  		radiometer_flags:SA\ overflow = "SAOVERFLOW" ;
  		radiometer_flags:Roughness\ correction\ failure = "ROUGH" ;
  		radiometer_flags:Solar\ flare\ contamination = "FLARE" ;
  		radiometer_flags:Pointing\ anomaly = "POINTING" ;
  		radiometer_flags:Tb\ consistency = "TBCONS" ;
  		radiometer_flags:Cold\ water = "COLDWATER" ;
  		radiometer_flags:RFI\ level = "TFTADIFF" ;
  		radiometer_flags:Moon/Galaxy\ contamination = "REFL_1STOKES" ;
  		radiometer_flags:RFI\ regional\ contamination = "RFI_REGION" ;
  		radiometer_flags:valid_min = 0U ;
  		radiometer_flags:valid_max = 0U ;
  	ubyte scat_rfi_flags(phony_dim_2, phony_dim_3, phony_dim_6) ;
  		scat_rfi_flags:long_name = "Scatterometer RFI flags" ;
  		scat_rfi_flags:valid_min = 0UB ;
  		scat_rfi_flags:valid_max = 0UB ;
  	uint scatterometer_flags(phony_dim_2, phony_dim_3) ;
  		scatterometer_flags:long_name = "Scatterometer data quality flags" ;
  		scatterometer_flags:valid_min = 0U ;
  		scatterometer_flags:valid_max = 0U ;
  		scatterometer_flags:RFI\ corruption\ of\ signal = "RFI" ;
  		scatterometer_flags:Rain\ in\ main\ beam = "RAIN" ;
  		scatterometer_flags:Negative\ TOA\ sigma0 = "NEGSIG" ;
  		scatterometer_flags:Non-nominal\ attitude = "BADATT" ;
  		scatterometer_flags:Faraday\ rotation\ removal = "FARADAY" ;
  } // group Aquarius\ Flags

group: Block\ Attributes {
  dimensions:
  	phony_dim_7 = 4083 ;
  	phony_dim_8 = 3 ;
  	phony_dim_9 = 4 ;
  variables:
  	ushort rad_samples(phony_dim_7, phony_dim_8, phony_dim_9) ;
  		rad_samples:long_name = "Number of radiometer samples per average" ;
  		rad_samples:valid_min = 0US ;
  		rad_samples:valid_max = 0US ;
  	ushort scat_samples(phony_dim_7, phony_dim_8) ;
  		scat_samples:long_name = "Number of scatterometer samples per average" ;
  		scat_samples:valid_min = 0US ;
  		scat_samples:valid_max = 0US ;
  	double sec(phony_dim_7) ;
  		sec:long_name = "Block time, seconds of day" ;
  		sec:valid_min = 0. ;
  		sec:valid_max = 0. ;
  		sec:units = "seconds" ;
  		sec:_FillValue = -9999. ;
  	double secGPS(phony_dim_7) ;
  		secGPS:long_name = "Block time, GPS time" ;
  		secGPS:valid_min = 0. ;
  		secGPS:valid_max = 0. ;
  		secGPS:units = "seconds" ;
  		secGPS:_FillValue = -9999. ;
  	float solar\ xray\ flux(phony_dim_7) ;
  		solar\ xray\ flux:long_name = "Solar xray flux (0.1 - 0.8 nanometers)" ;
  		solar\ xray\ flux:valid_min = 0.f ;
  		solar\ xray\ flux:valid_max = 0.f ;
  		solar\ xray\ flux:units = "watts/m2" ;
  		solar\ xray\ flux:_FillValue = -9999.f ;
  } // group Block\ Attributes

group: Converted\ Telemetry {
  dimensions:
  	phony_dim_10 = 4083 ;
  	phony_dim_11 = 85 ;
  	phony_dim_12 = 3 ;
  variables:
  	float rad_caltemps(phony_dim_10, phony_dim_11) ;
  		rad_caltemps:long_name = "Radiometer calibration temperatures" ;
  		rad_caltemps:valid_min = 0.f ;
  		rad_caltemps:valid_max = 0.f ;
  		rad_caltemps:_FillValue = -9999.f ;
  	float rad_ghh(phony_dim_10, phony_dim_12) ;
  		rad_ghh:long_name = "Radiometer HH gain" ;
  		rad_ghh:valid_min = 0.f ;
  		rad_ghh:valid_max = 0.f ;
  		rad_ghh:_FillValue = -9999.f ;
  	float rad_gmm(phony_dim_10, phony_dim_12) ;
  		rad_gmm:long_name = "Radiometer MM gain" ;
  		rad_gmm:valid_min = 0.f ;
  		rad_gmm:valid_max = 0.f ;
  		rad_gmm:_FillValue = -9999.f ;
  	float rad_gpp(phony_dim_10, phony_dim_12) ;
  		rad_gpp:long_name = "Radiometer PP gain" ;
  		rad_gpp:valid_min = 0.f ;
  		rad_gpp:valid_max = 0.f ;
  		rad_gpp:_FillValue = -9999.f ;
  	float rad_gvv(phony_dim_10, phony_dim_12) ;
  		rad_gvv:long_name = "Radiometer VV gain" ;
  		rad_gvv:valid_min = 0.f ;
  		rad_gvv:valid_max = 0.f ;
  		rad_gvv:_FillValue = -9999.f ;
  	float rad_oh(phony_dim_10, phony_dim_12) ;
  		rad_oh:long_name = "Radiometer H offset" ;
  		rad_oh:valid_min = 0.f ;
  		rad_oh:valid_max = 0.f ;
  		rad_oh:_FillValue = -9999.f ;
  	float rad_om(phony_dim_10, phony_dim_12) ;
  		rad_om:long_name = "Radiometer M offset" ;
  		rad_om:valid_min = 0.f ;
  		rad_om:valid_max = 0.f ;
  		rad_om:_FillValue = -9999.f ;
  	float rad_op(phony_dim_10, phony_dim_12) ;
  		rad_op:long_name = "Radiometer P offset" ;
  		rad_op:valid_max = 0.f ;
  		rad_op:_FillValue = -9999.f ;
  		rad_op:valid_min = 0.f ;
  	float rad_ov(phony_dim_10, phony_dim_12) ;
  		rad_ov:long_name = "Radiometer V offset" ;
  		rad_ov:valid_min = 0.f ;
  		rad_ov:valid_max = 0.f ;
  		rad_ov:_FillValue = -9999.f ;
  } // group Converted\ Telemetry

group: Navigation {
  dimensions:
  	phony_dim_13 = 4083 ;
  	phony_dim_14 = 3 ;
  	phony_dim_15 = 4 ;
  variables:
  	ubyte acs_mode(phony_dim_13) ;
  		acs_mode:long_name = "ACS Control Mode" ;
  		acs_mode:valid_min = 3UB ;
  		acs_mode:valid_max = 6UB ;
  	double att_ang(phony_dim_13, phony_dim_14) ;
  		att_ang:long_name = "Spacecraft roll, pitch, yaw" ;
  		att_ang:valid_min = -180. ;
  		att_ang:valid_max = 180. ;
  		att_ang:units = "degrees" ;
  		att_ang:_FillValue = -9999. ;
  	float beam_clat(phony_dim_13, phony_dim_14) ;
  		beam_clat:long_name = "Beam Center Latitude" ;
  		beam_clat:valid_min = -90.f ;
  		beam_clat:valid_max = 90.f ;
  		beam_clat:units = "degrees" ;
  		beam_clat:_FillValue = -9999.f ;
  	float beam_clon(phony_dim_13, phony_dim_14) ;
  		beam_clon:long_name = "Beam Center Longitude" ;
  		beam_clon:valid_min = -180.f ;
  		beam_clon:valid_max = 180.f ;
  		beam_clon:units = "degrees" ;
  		beam_clon:_FillValue = -9999.f ;
  	float cellatfoot(phony_dim_13, phony_dim_14, phony_dim_15) ;
  		cellatfoot:long_name = "Geodectic Latitudes (3 dB)" ;
  		cellatfoot:valid_min = -90.f ;
  		cellatfoot:valid_max = 90.f ;
  		cellatfoot:units = "degrees" ;
  		cellatfoot:_FillValue = -9999.f ;
  	float cellonfoot(phony_dim_13, phony_dim_14, phony_dim_15) ;
  		cellonfoot:long_name = "East Longitudes (3 dB)" ;
  		cellonfoot:valid_min = -180.f ;
  		cellonfoot:valid_max = 180.f ;
  		cellonfoot:units = "degrees" ;
  		cellonfoot:_FillValue = -9999.f ;
  	float celphi(phony_dim_13, phony_dim_14) ;
  		celphi:long_name = "Boresight Earth Azimuth Angle" ;
  		celphi:valid_min = -180.f ;
  		celphi:valid_max = 180.f ;
  		celphi:units = "degrees" ;
  		celphi:_FillValue = -9999.f ;
  	float celtht(phony_dim_13, phony_dim_14) ;
  		celtht:long_name = "Boresight Earth Incidence Angle" ;
  		celtht:valid_min = -180.f ;
  		celtht:valid_max = 180.f ;
  		celtht:units = "degrees" ;
  		celtht:_FillValue = -9999.f ;
  	float glxlat(phony_dim_13, phony_dim_14) ;
  		glxlat:long_name = "Galaxy Declination (J2000)" ;
  		glxlat:valid_min = -90.f ;
  		glxlat:valid_max = 90.f ;
  		glxlat:units = "degrees" ;
  		glxlat:_FillValue = -9999.f ;
  	float glxlon(phony_dim_13, phony_dim_14) ;
  		glxlon:long_name = "Galaxy Right Ascention (J2000)" ;
  		glxlon:valid_min = -180.f ;
  		glxlon:valid_max = 180.f ;
  		glxlon:units = "degrees" ;
  		glxlon:_FillValue = -9999.f ;
  	double moond(phony_dim_13, phony_dim_14) ;
  		moond:long_name = "Earth-to-Moon unit vector (eci)" ;
  		moond:valid_min = 0. ;
  		moond:valid_max = 0. ;
  		moond:_FillValue = -9999. ;
  	float moonglt(phony_dim_13, phony_dim_14) ;
  		moonglt:long_name = "Moon Glint Angle" ;
  		moonglt:valid_min = -180.f ;
  		moonglt:valid_max = 180.f ;
  		moonglt:units = "degrees" ;
  		moonglt:_FillValue = -9999.f ;
  	double orb_pos(phony_dim_13, phony_dim_14) ;
  		orb_pos:long_name = "Orbital position vector" ;
  		orb_pos:valid_min = -7100000. ;
  		orb_pos:valid_max = 7100000. ;
  		orb_pos:units = "meters" ;
  		orb_pos:_FillValue = -9999. ;
  	double orb_vel(phony_dim_13, phony_dim_14) ;
  		orb_vel:long_name = "Orbital velocity vector" ;
  		orb_vel:valid_min = -7600. ;
  		orb_vel:valid_max = 7600. ;
  		orb_vel:units = "meters per second" ;
  		orb_vel:_FillValue = -9999. ;
  	double scalt(phony_dim_13) ;
  		scalt:long_name = "Spacecraft altitude" ;
  		scalt:valid_min = 0. ;
  		scalt:valid_max = 0. ;
  		scalt:units = "meters" ;
  		scalt:_FillValue = -9999. ;
  	float scat_beam_clat(phony_dim_13, phony_dim_14) ;
  		scat_beam_clat:long_name = "Scatterometer Beam Center Latitude" ;
  		scat_beam_clat:valid_min = -90.f ;
  		scat_beam_clat:valid_max = 90.f ;
  		scat_beam_clat:units = "degrees" ;
  		scat_beam_clat:_FillValue = -9999.f ;
  	float scat_beam_clon(phony_dim_13, phony_dim_14) ;
  		scat_beam_clon:long_name = "Scatterometer Beam Center Longitude" ;
  		scat_beam_clon:valid_min = -180.f ;
  		scat_beam_clon:valid_max = 180.f ;
  		scat_beam_clon:units = "degrees" ;
  		scat_beam_clon:_FillValue = -9999.f ;
  	float scat_latfoot(phony_dim_13, phony_dim_14, phony_dim_15) ;
  		scat_latfoot:long_name = "Scatterometer Latitude Footprint" ;
  		scat_latfoot:valid_min = -90.f ;
  		scat_latfoot:valid_max = 90.f ;
  		scat_latfoot:units = "degrees" ;
  		scat_latfoot:_FillValue = -9999.f ;
  	float scat_lonfoot(phony_dim_13, phony_dim_14, phony_dim_15) ;
  		scat_lonfoot:long_name = "Scatterometer Longitude Footprint" ;
  		scat_lonfoot:valid_min = -180.f ;
  		scat_lonfoot:valid_max = 180.f ;
  		scat_lonfoot:units = "degrees" ;
  		scat_lonfoot:_FillValue = -9999.f ;
  	float scat_polarization_roll(phony_dim_13, phony_dim_14) ;
  		scat_polarization_roll:long_name = "Scatterometer Polarization Roll Angle" ;
  		scat_polarization_roll:valid_min = -180.f ;
  		scat_polarization_roll:valid_max = 180.f ;
  		scat_polarization_roll:units = "degrees" ;
  		scat_polarization_roll:_FillValue = -9999.f ;
  	double sclat(phony_dim_13) ;
  		sclat:long_name = "Spacecraft nadir point latitude" ;
  		sclat:valid_min = -90. ;
  		sclat:valid_max = 90. ;
  		sclat:units = "degrees" ;
  		sclat:_FillValue = -9999. ;
  	double sclon(phony_dim_13) ;
  		sclon:long_name = "Spacecraft nadir point longitude" ;
  		sclon:valid_min = -180. ;
  		sclon:valid_max = 180. ;
  		sclon:units = "degrees" ;
  		sclon:_FillValue = -9999. ;
  	double sund(phony_dim_13, phony_dim_14) ;
  		sund:long_name = "Earth-to-Sun unit vector (eci)" ;
  		sund:_FillValue = -9999. ;
  		sund:valid_min = 0. ;
  		sund:valid_max = 0. ;
  	float sunglt(phony_dim_13, phony_dim_14) ;
  		sunglt:long_name = "Sun Glint Angle" ;
  		sunglt:valid_min = -180.f ;
  		sunglt:valid_max = 180.f ;
  		sunglt:units = "degrees" ;
  		sunglt:_FillValue = -9999.f ;
  	float sunphi(phony_dim_13, phony_dim_14) ;
  		sunphi:long_name = "Sun Vector Earth Azimuth Angle" ;
  		sunphi:valid_min = -180.f ;
  		sunphi:valid_max = 180.f ;
  		sunphi:units = "degrees" ;
  		sunphi:_FillValue = -9999.f ;
  	double sunr(phony_dim_13, phony_dim_14) ;
  		sunr:long_name = "Sun reflection unit vector (eci)" ;
  		sunr:valid_min = 0. ;
  		sunr:valid_max = 0. ;
  		sunr:_FillValue = -9999. ;
  	float suntht(phony_dim_13, phony_dim_14) ;
  		suntht:long_name = "Sun Vector Earth Incidence Angle" ;
  		suntht:valid_min = -180.f ;
  		suntht:valid_max = 180.f ;
  		suntht:units = "degrees" ;
  		suntht:_FillValue = -9999.f ;
  	double zang(phony_dim_13) ;
  		zang:long_name = "Intra-Orbit Angle" ;
  		zang:valid_min = -180. ;
  		zang:valid_max = 180. ;
  		zang:units = "degrees" ;
  		zang:_FillValue = -9999. ;
  } // group Navigation
}
