// -*-C++-*-

// Purpose: CDL file to demonstrate best practices for rectangular gridded datasets
// Part of an ongoing project by NASA's Dataset Interoperability Working Group (DIWG)
// Comments, questions, suggestions to fxm

// Usage:
// ncgen             -b -o global_rectangular.nc global_rectangular.cdl # netCDF3
// ncgen -k netCDF-4 -b -o global_rectangular.nc global_rectangular.cdl # netCDF4

// URL: 
// git clone http://github.com/diwg/diwg.git
// http://github.com/diwg/diwg/global_rectangular.cdl

netcdf global_rectangular {
 dimensions:
  longitude = 2 ;
  latitude = 2 ;
  time = UNLIMITED ; // time = 1 for files w/one time slice
  
 variables:
  // Grid coordinates are double precision to retain accuracy during remapping
  double longitude(longitude);
  longitude:standard_name = "longitude";
  longitude:units = "degrees_east";
  longitude:axis = "X";

  double latitude(latitude) ;
  latitude:standard_name = "latitude";
  latitude:units = "degrees_north";  
  latitude:axis = "Y";

  short TB(time, latitude, longitude);
 TB:long_name = "brightness temperature";
 TB:standard_name = "brightness_temperature";
 TB:units = "kelvin";
 TB:scale_factor = 0.01f;
 TB:add_offset = 0.0f;
 TB:packing_convention = "netCDF";
 TB:packing_convention_description = "unpacked = scale_factor*packed + add_offset";
 TB:grid_mapping = "crs";
  
  byte TB_num_samples(time, latitude, longitude);
 TB_num_samples:long_name = "brightness temperature number of samples";
 TB_num_samples:units = "1";
 TB_num_samples:grid_mapping = "crs";

  char crs ;
  // CF Grid Mappings: http://cfconventions.org/Data/cf-conventions/cf-conventions-1.7/build/apf.html
  // fxm: Projection data is meaningless for global gridded data (move to a different template file)
 crs:grid_mapping_name = "lambert_cylindrical_equal_area" ;
 crs:crs_wkt = "PROJCS[
	    BASE_GEODGCS[\"WGS 84\",
	        DATUM[ \"World Geodetic System 1984\",
		    ELLIPSOID[\"WGS 84\",
		    6378137,298.257223563,
		    LENGTHUNIT[\"metre\",\"1.0\"]]]],
    	    ID[\"EPSG,6933\"]]" ;

 data:
  longitude=0.,360.;
  latitude=-90.,90.;
  TB=1,2,3,4;
  TB_num_samples='1','2','3','4';
} // end netcdf
